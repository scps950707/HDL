
module pipealu_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [33:0] carry;
  wire   [32:0] B_AS;
  assign carry[0] = ADD_SUB;

  FADDX1 U1_31 ( .A(A[31]), .B(B_AS[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B_AS[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B_AS[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B_AS[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B_AS[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B_AS[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B_AS[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B_AS[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B_AS[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B_AS[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B_AS[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B_AS[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B_AS[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B_AS[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B_AS[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B_AS[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B_AS[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FADDX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FADDX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FADDX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FADDX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FADDX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FADDX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FADDX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FADDX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0]) );
  XOR2X1 U1 ( .IN1(carry[0]), .IN2(carry[32]), .Q(SUM[32]) );
  XOR2X1 U2 ( .IN1(B[9]), .IN2(carry[0]), .Q(B_AS[9]) );
  XOR2X1 U3 ( .IN1(B[8]), .IN2(carry[0]), .Q(B_AS[8]) );
  XOR2X1 U4 ( .IN1(B[7]), .IN2(carry[0]), .Q(B_AS[7]) );
  XOR2X1 U5 ( .IN1(B[6]), .IN2(carry[0]), .Q(B_AS[6]) );
  XOR2X1 U6 ( .IN1(B[5]), .IN2(carry[0]), .Q(B_AS[5]) );
  XOR2X1 U7 ( .IN1(B[4]), .IN2(carry[0]), .Q(B_AS[4]) );
  XOR2X1 U8 ( .IN1(B[3]), .IN2(carry[0]), .Q(B_AS[3]) );
  XOR2X1 U9 ( .IN1(B[31]), .IN2(carry[0]), .Q(B_AS[31]) );
  XOR2X1 U10 ( .IN1(B[30]), .IN2(carry[0]), .Q(B_AS[30]) );
  XOR2X1 U11 ( .IN1(B[2]), .IN2(carry[0]), .Q(B_AS[2]) );
  XOR2X1 U12 ( .IN1(B[29]), .IN2(carry[0]), .Q(B_AS[29]) );
  XOR2X1 U13 ( .IN1(B[28]), .IN2(carry[0]), .Q(B_AS[28]) );
  XOR2X1 U14 ( .IN1(B[27]), .IN2(carry[0]), .Q(B_AS[27]) );
  XOR2X1 U15 ( .IN1(B[26]), .IN2(carry[0]), .Q(B_AS[26]) );
  XOR2X1 U16 ( .IN1(B[25]), .IN2(carry[0]), .Q(B_AS[25]) );
  XOR2X1 U17 ( .IN1(B[24]), .IN2(carry[0]), .Q(B_AS[24]) );
  XOR2X1 U18 ( .IN1(B[23]), .IN2(carry[0]), .Q(B_AS[23]) );
  XOR2X1 U19 ( .IN1(B[22]), .IN2(carry[0]), .Q(B_AS[22]) );
  XOR2X1 U20 ( .IN1(B[21]), .IN2(carry[0]), .Q(B_AS[21]) );
  XOR2X1 U21 ( .IN1(B[20]), .IN2(carry[0]), .Q(B_AS[20]) );
  XOR2X1 U22 ( .IN1(B[1]), .IN2(carry[0]), .Q(B_AS[1]) );
  XOR2X1 U23 ( .IN1(B[19]), .IN2(carry[0]), .Q(B_AS[19]) );
  XOR2X1 U24 ( .IN1(B[18]), .IN2(carry[0]), .Q(B_AS[18]) );
  XOR2X1 U25 ( .IN1(B[17]), .IN2(carry[0]), .Q(B_AS[17]) );
  XOR2X1 U26 ( .IN1(B[16]), .IN2(carry[0]), .Q(B_AS[16]) );
  XOR2X1 U27 ( .IN1(B[15]), .IN2(carry[0]), .Q(B_AS[15]) );
  XOR2X1 U28 ( .IN1(B[14]), .IN2(carry[0]), .Q(B_AS[14]) );
  XOR2X1 U29 ( .IN1(B[13]), .IN2(carry[0]), .Q(B_AS[13]) );
  XOR2X1 U30 ( .IN1(B[12]), .IN2(carry[0]), .Q(B_AS[12]) );
  XOR2X1 U31 ( .IN1(B[11]), .IN2(carry[0]), .Q(B_AS[11]) );
  XOR2X1 U32 ( .IN1(B[10]), .IN2(carry[0]), .Q(B_AS[10]) );
  XOR2X1 U33 ( .IN1(B[0]), .IN2(carry[0]), .Q(B_AS[0]) );
endmodule


module pipealu ( instr, AluOut, Zero, clk, Carryout, Overflow, rst );
  input [15:0] instr;
  output [31:0] AluOut;
  input clk, rst;
  output Zero, Carryout, Overflow;
  wire   N15, N16, N17, N18, N19, N20, N21, N22, \regfile[15][31] ,
         \regfile[15][30] , \regfile[15][29] , \regfile[15][28] ,
         \regfile[15][27] , \regfile[15][26] , \regfile[15][25] ,
         \regfile[15][24] , \regfile[15][23] , \regfile[15][22] ,
         \regfile[15][21] , \regfile[15][20] , \regfile[15][19] ,
         \regfile[15][18] , \regfile[15][17] , \regfile[15][16] ,
         \regfile[15][15] , \regfile[15][14] , \regfile[15][13] ,
         \regfile[15][12] , \regfile[15][11] , \regfile[15][10] ,
         \regfile[15][9] , \regfile[15][8] , \regfile[15][7] ,
         \regfile[15][6] , \regfile[15][5] , \regfile[15][4] ,
         \regfile[15][3] , \regfile[15][2] , \regfile[15][1] ,
         \regfile[15][0] , \regfile[14][31] , \regfile[14][30] ,
         \regfile[14][29] , \regfile[14][28] , \regfile[14][27] ,
         \regfile[14][26] , \regfile[14][25] , \regfile[14][24] ,
         \regfile[14][23] , \regfile[14][22] , \regfile[14][21] ,
         \regfile[14][20] , \regfile[14][19] , \regfile[14][18] ,
         \regfile[14][17] , \regfile[14][16] , \regfile[14][15] ,
         \regfile[14][14] , \regfile[14][13] , \regfile[14][12] ,
         \regfile[14][11] , \regfile[14][10] , \regfile[14][9] ,
         \regfile[14][8] , \regfile[14][7] , \regfile[14][6] ,
         \regfile[14][5] , \regfile[14][4] , \regfile[14][3] ,
         \regfile[14][2] , \regfile[14][1] , \regfile[14][0] ,
         \regfile[13][31] , \regfile[13][30] , \regfile[13][29] ,
         \regfile[13][28] , \regfile[13][27] , \regfile[13][26] ,
         \regfile[13][25] , \regfile[13][24] , \regfile[13][23] ,
         \regfile[13][22] , \regfile[13][21] , \regfile[13][20] ,
         \regfile[13][19] , \regfile[13][18] , \regfile[13][17] ,
         \regfile[13][16] , \regfile[13][15] , \regfile[13][14] ,
         \regfile[13][13] , \regfile[13][12] , \regfile[13][11] ,
         \regfile[13][10] , \regfile[13][9] , \regfile[13][8] ,
         \regfile[13][7] , \regfile[13][6] , \regfile[13][5] ,
         \regfile[13][4] , \regfile[13][3] , \regfile[13][2] ,
         \regfile[13][1] , \regfile[13][0] , \regfile[12][31] ,
         \regfile[12][30] , \regfile[12][29] , \regfile[12][28] ,
         \regfile[12][27] , \regfile[12][26] , \regfile[12][25] ,
         \regfile[12][24] , \regfile[12][23] , \regfile[12][22] ,
         \regfile[12][21] , \regfile[12][20] , \regfile[12][19] ,
         \regfile[12][18] , \regfile[12][17] , \regfile[12][16] ,
         \regfile[12][15] , \regfile[12][14] , \regfile[12][13] ,
         \regfile[12][12] , \regfile[12][11] , \regfile[12][10] ,
         \regfile[12][9] , \regfile[12][8] , \regfile[12][7] ,
         \regfile[12][6] , \regfile[12][5] , \regfile[12][4] ,
         \regfile[12][3] , \regfile[12][2] , \regfile[12][1] ,
         \regfile[12][0] , \regfile[11][31] , \regfile[11][30] ,
         \regfile[11][29] , \regfile[11][28] , \regfile[11][27] ,
         \regfile[11][26] , \regfile[11][25] , \regfile[11][24] ,
         \regfile[11][23] , \regfile[11][22] , \regfile[11][21] ,
         \regfile[11][20] , \regfile[11][19] , \regfile[11][18] ,
         \regfile[11][17] , \regfile[11][16] , \regfile[11][15] ,
         \regfile[11][14] , \regfile[11][13] , \regfile[11][12] ,
         \regfile[11][11] , \regfile[11][10] , \regfile[11][9] ,
         \regfile[11][8] , \regfile[11][7] , \regfile[11][6] ,
         \regfile[11][5] , \regfile[11][4] , \regfile[11][3] ,
         \regfile[11][2] , \regfile[11][1] , \regfile[11][0] ,
         \regfile[10][31] , \regfile[10][30] , \regfile[10][29] ,
         \regfile[10][28] , \regfile[10][27] , \regfile[10][26] ,
         \regfile[10][25] , \regfile[10][24] , \regfile[10][23] ,
         \regfile[10][22] , \regfile[10][21] , \regfile[10][20] ,
         \regfile[10][19] , \regfile[10][18] , \regfile[10][17] ,
         \regfile[10][16] , \regfile[10][15] , \regfile[10][14] ,
         \regfile[10][13] , \regfile[10][12] , \regfile[10][11] ,
         \regfile[10][10] , \regfile[10][9] , \regfile[10][8] ,
         \regfile[10][7] , \regfile[10][6] , \regfile[10][5] ,
         \regfile[10][4] , \regfile[10][3] , \regfile[10][2] ,
         \regfile[10][1] , \regfile[10][0] , \regfile[9][31] ,
         \regfile[9][30] , \regfile[9][29] , \regfile[9][28] ,
         \regfile[9][27] , \regfile[9][26] , \regfile[9][25] ,
         \regfile[9][24] , \regfile[9][23] , \regfile[9][22] ,
         \regfile[9][21] , \regfile[9][20] , \regfile[9][19] ,
         \regfile[9][18] , \regfile[9][17] , \regfile[9][16] ,
         \regfile[9][15] , \regfile[9][14] , \regfile[9][13] ,
         \regfile[9][12] , \regfile[9][11] , \regfile[9][10] , \regfile[9][9] ,
         \regfile[9][8] , \regfile[9][7] , \regfile[9][6] , \regfile[9][5] ,
         \regfile[9][4] , \regfile[9][3] , \regfile[9][2] , \regfile[9][1] ,
         \regfile[9][0] , \regfile[8][31] , \regfile[8][30] , \regfile[8][29] ,
         \regfile[8][28] , \regfile[8][27] , \regfile[8][26] ,
         \regfile[8][25] , \regfile[8][24] , \regfile[8][23] ,
         \regfile[8][22] , \regfile[8][21] , \regfile[8][20] ,
         \regfile[8][19] , \regfile[8][18] , \regfile[8][17] ,
         \regfile[8][16] , \regfile[8][15] , \regfile[8][14] ,
         \regfile[8][13] , \regfile[8][12] , \regfile[8][11] ,
         \regfile[8][10] , \regfile[8][9] , \regfile[8][8] , \regfile[8][7] ,
         \regfile[8][6] , \regfile[8][5] , \regfile[8][4] , \regfile[8][3] ,
         \regfile[8][2] , \regfile[8][1] , \regfile[8][0] , \regfile[7][31] ,
         \regfile[7][30] , \regfile[7][29] , \regfile[7][28] ,
         \regfile[7][27] , \regfile[7][26] , \regfile[7][25] ,
         \regfile[7][24] , \regfile[7][23] , \regfile[7][22] ,
         \regfile[7][21] , \regfile[7][20] , \regfile[7][19] ,
         \regfile[7][18] , \regfile[7][17] , \regfile[7][16] ,
         \regfile[7][15] , \regfile[7][14] , \regfile[7][13] ,
         \regfile[7][12] , \regfile[7][11] , \regfile[7][10] , \regfile[7][9] ,
         \regfile[7][8] , \regfile[7][7] , \regfile[7][6] , \regfile[7][5] ,
         \regfile[7][4] , \regfile[7][3] , \regfile[7][2] , \regfile[7][1] ,
         \regfile[7][0] , \regfile[6][31] , \regfile[6][30] , \regfile[6][29] ,
         \regfile[6][28] , \regfile[6][27] , \regfile[6][26] ,
         \regfile[6][25] , \regfile[6][24] , \regfile[6][23] ,
         \regfile[6][22] , \regfile[6][21] , \regfile[6][20] ,
         \regfile[6][19] , \regfile[6][18] , \regfile[6][17] ,
         \regfile[6][16] , \regfile[6][15] , \regfile[6][14] ,
         \regfile[6][13] , \regfile[6][12] , \regfile[6][11] ,
         \regfile[6][10] , \regfile[6][9] , \regfile[6][8] , \regfile[6][7] ,
         \regfile[6][6] , \regfile[6][5] , \regfile[6][4] , \regfile[6][3] ,
         \regfile[6][2] , \regfile[6][1] , \regfile[6][0] , \regfile[5][31] ,
         \regfile[5][30] , \regfile[5][29] , \regfile[5][28] ,
         \regfile[5][27] , \regfile[5][26] , \regfile[5][25] ,
         \regfile[5][24] , \regfile[5][23] , \regfile[5][22] ,
         \regfile[5][21] , \regfile[5][20] , \regfile[5][19] ,
         \regfile[5][18] , \regfile[5][17] , \regfile[5][16] ,
         \regfile[5][15] , \regfile[5][14] , \regfile[5][13] ,
         \regfile[5][12] , \regfile[5][11] , \regfile[5][10] , \regfile[5][9] ,
         \regfile[5][8] , \regfile[5][7] , \regfile[5][6] , \regfile[5][5] ,
         \regfile[5][4] , \regfile[5][3] , \regfile[5][2] , \regfile[5][1] ,
         \regfile[5][0] , \regfile[4][31] , \regfile[4][30] , \regfile[4][29] ,
         \regfile[4][28] , \regfile[4][27] , \regfile[4][26] ,
         \regfile[4][25] , \regfile[4][24] , \regfile[4][23] ,
         \regfile[4][22] , \regfile[4][21] , \regfile[4][20] ,
         \regfile[4][19] , \regfile[4][18] , \regfile[4][17] ,
         \regfile[4][16] , \regfile[4][15] , \regfile[4][14] ,
         \regfile[4][13] , \regfile[4][12] , \regfile[4][11] ,
         \regfile[4][10] , \regfile[4][9] , \regfile[4][8] , \regfile[4][7] ,
         \regfile[4][6] , \regfile[4][5] , \regfile[4][4] , \regfile[4][3] ,
         \regfile[4][2] , \regfile[4][1] , \regfile[4][0] , \regfile[3][31] ,
         \regfile[3][30] , \regfile[3][29] , \regfile[3][28] ,
         \regfile[3][27] , \regfile[3][26] , \regfile[3][25] ,
         \regfile[3][24] , \regfile[3][23] , \regfile[3][22] ,
         \regfile[3][21] , \regfile[3][20] , \regfile[3][19] ,
         \regfile[3][18] , \regfile[3][17] , \regfile[3][16] ,
         \regfile[3][15] , \regfile[3][14] , \regfile[3][13] ,
         \regfile[3][12] , \regfile[3][11] , \regfile[3][10] , \regfile[3][9] ,
         \regfile[3][8] , \regfile[3][7] , \regfile[3][6] , \regfile[3][5] ,
         \regfile[3][4] , \regfile[3][3] , \regfile[3][2] , \regfile[3][1] ,
         \regfile[3][0] , \regfile[2][31] , \regfile[2][30] , \regfile[2][29] ,
         \regfile[2][28] , \regfile[2][27] , \regfile[2][26] ,
         \regfile[2][25] , \regfile[2][24] , \regfile[2][23] ,
         \regfile[2][22] , \regfile[2][21] , \regfile[2][20] ,
         \regfile[2][19] , \regfile[2][18] , \regfile[2][17] ,
         \regfile[2][16] , \regfile[2][15] , \regfile[2][14] ,
         \regfile[2][13] , \regfile[2][12] , \regfile[2][11] ,
         \regfile[2][10] , \regfile[2][9] , \regfile[2][8] , \regfile[2][7] ,
         \regfile[2][6] , \regfile[2][5] , \regfile[2][4] , \regfile[2][3] ,
         \regfile[2][2] , \regfile[2][1] , \regfile[2][0] , \regfile[1][31] ,
         \regfile[1][30] , \regfile[1][29] , \regfile[1][28] ,
         \regfile[1][27] , \regfile[1][26] , \regfile[1][25] ,
         \regfile[1][24] , \regfile[1][23] , \regfile[1][22] ,
         \regfile[1][21] , \regfile[1][20] , \regfile[1][19] ,
         \regfile[1][18] , \regfile[1][17] , \regfile[1][16] ,
         \regfile[1][15] , \regfile[1][14] , \regfile[1][13] ,
         \regfile[1][12] , \regfile[1][11] , \regfile[1][10] , \regfile[1][9] ,
         \regfile[1][8] , \regfile[1][7] , \regfile[1][6] , \regfile[1][5] ,
         \regfile[1][4] , \regfile[1][3] , \regfile[1][2] , \regfile[1][1] ,
         \regfile[1][0] , \regfile[0][31] , \regfile[0][30] , \regfile[0][29] ,
         \regfile[0][28] , \regfile[0][27] , \regfile[0][26] ,
         \regfile[0][25] , \regfile[0][24] , \regfile[0][23] ,
         \regfile[0][22] , \regfile[0][21] , \regfile[0][20] ,
         \regfile[0][19] , \regfile[0][18] , \regfile[0][17] ,
         \regfile[0][16] , \regfile[0][15] , \regfile[0][14] ,
         \regfile[0][13] , \regfile[0][12] , \regfile[0][11] ,
         \regfile[0][10] , \regfile[0][9] , \regfile[0][8] , \regfile[0][7] ,
         \regfile[0][6] , \regfile[0][5] , \regfile[0][4] , \regfile[0][3] ,
         \regfile[0][2] , \regfile[0][1] , \regfile[0][0] , N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N257, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318;
  wire   [31:0] IFID_A;
  wire   [31:0] IFID_B;
  assign N15 = instr[8];
  assign N16 = instr[9];
  assign N17 = instr[10];
  assign N18 = instr[11];
  assign N19 = instr[4];
  assign N20 = instr[5];
  assign N21 = instr[6];
  assign N22 = instr[7];

  DFFX1 Carryout_reg ( .D(n1317), .CLK(clk), .Q(Carryout) );
  DFFX1 \EX_dest_reg[3]  ( .D(instr[3]), .CLK(clk), .Q(n1315) );
  DFFX1 \EX_dest_reg[2]  ( .D(instr[2]), .CLK(clk), .Q(n1313) );
  DFFX1 \EX_dest_reg[1]  ( .D(instr[1]), .CLK(clk), .Q(n1316), .QN(n799) );
  DFFX1 \EX_dest_reg[0]  ( .D(instr[0]), .CLK(clk), .Q(n1314), .QN(n800) );
  DFFX1 Overflow_reg ( .D(N257), .CLK(clk), .Q(Overflow) );
  DFFX1 \AluOut_reg[31]  ( .D(n795), .CLK(clk), .Q(AluOut[31]), .QN(n251) );
  DFFARX1 \regfile_reg[0][31]  ( .D(n794), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][31] ) );
  DFFARX1 \regfile_reg[1][31]  ( .D(n793), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][31] ) );
  DFFARX1 \regfile_reg[2][31]  ( .D(n792), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][31] ) );
  DFFARX1 \regfile_reg[3][31]  ( .D(n791), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][31] ) );
  DFFARX1 \regfile_reg[4][31]  ( .D(n790), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][31] ) );
  DFFARX1 \regfile_reg[5][31]  ( .D(n789), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][31] ) );
  DFFARX1 \regfile_reg[6][31]  ( .D(n788), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][31] ) );
  DFFARX1 \regfile_reg[7][31]  ( .D(n787), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][31] ) );
  DFFARX1 \regfile_reg[8][31]  ( .D(n786), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][31] ) );
  DFFARX1 \regfile_reg[9][31]  ( .D(n785), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][31] ) );
  DFFARX1 \regfile_reg[10][31]  ( .D(n784), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][31] ) );
  DFFARX1 \regfile_reg[11][31]  ( .D(n783), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][31] ) );
  DFFARX1 \regfile_reg[12][31]  ( .D(n782), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][31] ) );
  DFFARX1 \regfile_reg[13][31]  ( .D(n781), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][31] ) );
  DFFARX1 \regfile_reg[14][31]  ( .D(n780), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][31] ) );
  DFFARX1 \regfile_reg[15][31]  ( .D(n779), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][31] ) );
  DFFX1 \AluOut_reg[30]  ( .D(n778), .CLK(clk), .Q(AluOut[30]), .QN(n246) );
  DFFARX1 \regfile_reg[0][30]  ( .D(n777), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][30] ) );
  DFFARX1 \regfile_reg[1][30]  ( .D(n776), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][30] ) );
  DFFARX1 \regfile_reg[2][30]  ( .D(n775), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][30] ) );
  DFFARX1 \regfile_reg[3][30]  ( .D(n774), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][30] ) );
  DFFARX1 \regfile_reg[4][30]  ( .D(n773), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][30] ) );
  DFFARX1 \regfile_reg[5][30]  ( .D(n772), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][30] ) );
  DFFARX1 \regfile_reg[6][30]  ( .D(n771), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][30] ) );
  DFFARX1 \regfile_reg[7][30]  ( .D(n770), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][30] ) );
  DFFARX1 \regfile_reg[8][30]  ( .D(n769), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][30] ) );
  DFFARX1 \regfile_reg[9][30]  ( .D(n768), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][30] ) );
  DFFARX1 \regfile_reg[10][30]  ( .D(n767), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][30] ) );
  DFFARX1 \regfile_reg[11][30]  ( .D(n766), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][30] ) );
  DFFARX1 \regfile_reg[12][30]  ( .D(n765), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][30] ) );
  DFFARX1 \regfile_reg[13][30]  ( .D(n764), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][30] ) );
  DFFARX1 \regfile_reg[14][30]  ( .D(n763), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][30] ) );
  DFFARX1 \regfile_reg[15][30]  ( .D(n762), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][30] ) );
  DFFX1 \AluOut_reg[29]  ( .D(n761), .CLK(clk), .Q(AluOut[29]), .QN(n245) );
  DFFARX1 \regfile_reg[0][29]  ( .D(n760), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][29] ) );
  DFFARX1 \regfile_reg[1][29]  ( .D(n759), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][29] ) );
  DFFARX1 \regfile_reg[2][29]  ( .D(n758), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][29] ) );
  DFFARX1 \regfile_reg[3][29]  ( .D(n757), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][29] ) );
  DFFARX1 \regfile_reg[4][29]  ( .D(n756), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][29] ) );
  DFFARX1 \regfile_reg[5][29]  ( .D(n755), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][29] ) );
  DFFARX1 \regfile_reg[6][29]  ( .D(n754), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][29] ) );
  DFFARX1 \regfile_reg[7][29]  ( .D(n753), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][29] ) );
  DFFARX1 \regfile_reg[8][29]  ( .D(n752), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][29] ) );
  DFFARX1 \regfile_reg[9][29]  ( .D(n751), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][29] ) );
  DFFARX1 \regfile_reg[10][29]  ( .D(n750), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][29] ) );
  DFFARX1 \regfile_reg[11][29]  ( .D(n749), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][29] ) );
  DFFARX1 \regfile_reg[12][29]  ( .D(n748), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][29] ) );
  DFFARX1 \regfile_reg[13][29]  ( .D(n747), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][29] ) );
  DFFARX1 \regfile_reg[14][29]  ( .D(n746), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][29] ) );
  DFFARX1 \regfile_reg[15][29]  ( .D(n745), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][29] ) );
  DFFX1 \AluOut_reg[28]  ( .D(n744), .CLK(clk), .Q(AluOut[28]), .QN(n244) );
  DFFARX1 \regfile_reg[0][28]  ( .D(n743), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][28] ) );
  DFFARX1 \regfile_reg[1][28]  ( .D(n742), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][28] ) );
  DFFARX1 \regfile_reg[2][28]  ( .D(n741), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][28] ) );
  DFFARX1 \regfile_reg[3][28]  ( .D(n740), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][28] ) );
  DFFARX1 \regfile_reg[4][28]  ( .D(n739), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][28] ) );
  DFFARX1 \regfile_reg[5][28]  ( .D(n738), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][28] ) );
  DFFARX1 \regfile_reg[6][28]  ( .D(n737), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][28] ) );
  DFFARX1 \regfile_reg[7][28]  ( .D(n736), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][28] ) );
  DFFARX1 \regfile_reg[8][28]  ( .D(n735), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][28] ) );
  DFFARX1 \regfile_reg[9][28]  ( .D(n734), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][28] ) );
  DFFARX1 \regfile_reg[10][28]  ( .D(n733), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][28] ) );
  DFFARX1 \regfile_reg[11][28]  ( .D(n732), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][28] ) );
  DFFARX1 \regfile_reg[12][28]  ( .D(n731), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][28] ) );
  DFFARX1 \regfile_reg[13][28]  ( .D(n730), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][28] ) );
  DFFARX1 \regfile_reg[14][28]  ( .D(n729), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][28] ) );
  DFFARX1 \regfile_reg[15][28]  ( .D(n728), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][28] ) );
  DFFX1 \AluOut_reg[27]  ( .D(n727), .CLK(clk), .Q(AluOut[27]), .QN(n243) );
  DFFARX1 \regfile_reg[0][27]  ( .D(n726), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][27] ) );
  DFFARX1 \regfile_reg[1][27]  ( .D(n725), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][27] ) );
  DFFARX1 \regfile_reg[2][27]  ( .D(n724), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][27] ) );
  DFFARX1 \regfile_reg[3][27]  ( .D(n723), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][27] ) );
  DFFARX1 \regfile_reg[4][27]  ( .D(n722), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][27] ) );
  DFFARX1 \regfile_reg[5][27]  ( .D(n721), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][27] ) );
  DFFARX1 \regfile_reg[6][27]  ( .D(n720), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][27] ) );
  DFFARX1 \regfile_reg[7][27]  ( .D(n719), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][27] ) );
  DFFARX1 \regfile_reg[8][27]  ( .D(n718), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][27] ) );
  DFFARX1 \regfile_reg[9][27]  ( .D(n717), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][27] ) );
  DFFARX1 \regfile_reg[10][27]  ( .D(n716), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][27] ) );
  DFFARX1 \regfile_reg[11][27]  ( .D(n715), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][27] ) );
  DFFARX1 \regfile_reg[12][27]  ( .D(n714), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][27] ) );
  DFFARX1 \regfile_reg[13][27]  ( .D(n713), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][27] ) );
  DFFARX1 \regfile_reg[14][27]  ( .D(n712), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][27] ) );
  DFFARX1 \regfile_reg[15][27]  ( .D(n711), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][27] ) );
  DFFX1 \AluOut_reg[26]  ( .D(n710), .CLK(clk), .Q(AluOut[26]), .QN(n242) );
  DFFARX1 \regfile_reg[0][26]  ( .D(n709), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][26] ) );
  DFFARX1 \regfile_reg[1][26]  ( .D(n708), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][26] ) );
  DFFARX1 \regfile_reg[2][26]  ( .D(n707), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][26] ) );
  DFFARX1 \regfile_reg[3][26]  ( .D(n706), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][26] ) );
  DFFARX1 \regfile_reg[4][26]  ( .D(n705), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][26] ) );
  DFFARX1 \regfile_reg[5][26]  ( .D(n704), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][26] ) );
  DFFARX1 \regfile_reg[6][26]  ( .D(n703), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][26] ) );
  DFFARX1 \regfile_reg[7][26]  ( .D(n702), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][26] ) );
  DFFARX1 \regfile_reg[8][26]  ( .D(n701), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][26] ) );
  DFFARX1 \regfile_reg[9][26]  ( .D(n700), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][26] ) );
  DFFARX1 \regfile_reg[10][26]  ( .D(n699), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][26] ) );
  DFFARX1 \regfile_reg[11][26]  ( .D(n698), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][26] ) );
  DFFARX1 \regfile_reg[12][26]  ( .D(n697), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][26] ) );
  DFFARX1 \regfile_reg[13][26]  ( .D(n696), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][26] ) );
  DFFARX1 \regfile_reg[14][26]  ( .D(n695), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][26] ) );
  DFFARX1 \regfile_reg[15][26]  ( .D(n694), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][26] ) );
  DFFX1 \AluOut_reg[25]  ( .D(n693), .CLK(clk), .Q(AluOut[25]), .QN(n241) );
  DFFARX1 \regfile_reg[0][25]  ( .D(n692), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][25] ) );
  DFFARX1 \regfile_reg[1][25]  ( .D(n691), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][25] ) );
  DFFARX1 \regfile_reg[2][25]  ( .D(n690), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][25] ) );
  DFFARX1 \regfile_reg[3][25]  ( .D(n689), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][25] ) );
  DFFARX1 \regfile_reg[4][25]  ( .D(n688), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][25] ) );
  DFFARX1 \regfile_reg[5][25]  ( .D(n687), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][25] ) );
  DFFARX1 \regfile_reg[6][25]  ( .D(n686), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][25] ) );
  DFFARX1 \regfile_reg[7][25]  ( .D(n685), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][25] ) );
  DFFARX1 \regfile_reg[8][25]  ( .D(n684), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][25] ) );
  DFFARX1 \regfile_reg[9][25]  ( .D(n683), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][25] ) );
  DFFARX1 \regfile_reg[10][25]  ( .D(n682), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][25] ) );
  DFFARX1 \regfile_reg[11][25]  ( .D(n681), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][25] ) );
  DFFARX1 \regfile_reg[12][25]  ( .D(n680), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][25] ) );
  DFFARX1 \regfile_reg[13][25]  ( .D(n679), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][25] ) );
  DFFARX1 \regfile_reg[14][25]  ( .D(n678), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][25] ) );
  DFFARX1 \regfile_reg[15][25]  ( .D(n677), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][25] ) );
  DFFX1 \AluOut_reg[24]  ( .D(n676), .CLK(clk), .Q(AluOut[24]), .QN(n240) );
  DFFARX1 \regfile_reg[0][24]  ( .D(n675), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][24] ) );
  DFFARX1 \regfile_reg[1][24]  ( .D(n674), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][24] ) );
  DFFARX1 \regfile_reg[2][24]  ( .D(n673), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][24] ) );
  DFFARX1 \regfile_reg[3][24]  ( .D(n672), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][24] ) );
  DFFARX1 \regfile_reg[4][24]  ( .D(n671), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][24] ) );
  DFFARX1 \regfile_reg[5][24]  ( .D(n670), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][24] ) );
  DFFARX1 \regfile_reg[6][24]  ( .D(n669), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][24] ) );
  DFFARX1 \regfile_reg[7][24]  ( .D(n668), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][24] ) );
  DFFARX1 \regfile_reg[8][24]  ( .D(n667), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][24] ) );
  DFFARX1 \regfile_reg[9][24]  ( .D(n666), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][24] ) );
  DFFARX1 \regfile_reg[10][24]  ( .D(n665), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][24] ) );
  DFFARX1 \regfile_reg[11][24]  ( .D(n664), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][24] ) );
  DFFARX1 \regfile_reg[12][24]  ( .D(n663), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][24] ) );
  DFFARX1 \regfile_reg[13][24]  ( .D(n662), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][24] ) );
  DFFARX1 \regfile_reg[14][24]  ( .D(n661), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][24] ) );
  DFFARX1 \regfile_reg[15][24]  ( .D(n660), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][24] ) );
  DFFX1 \AluOut_reg[23]  ( .D(n659), .CLK(clk), .Q(AluOut[23]), .QN(n239) );
  DFFARX1 \regfile_reg[0][23]  ( .D(n658), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][23] ) );
  DFFARX1 \regfile_reg[1][23]  ( .D(n657), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][23] ) );
  DFFARX1 \regfile_reg[2][23]  ( .D(n656), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][23] ) );
  DFFARX1 \regfile_reg[3][23]  ( .D(n655), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][23] ) );
  DFFARX1 \regfile_reg[4][23]  ( .D(n654), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][23] ) );
  DFFARX1 \regfile_reg[5][23]  ( .D(n653), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][23] ) );
  DFFARX1 \regfile_reg[6][23]  ( .D(n652), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][23] ) );
  DFFARX1 \regfile_reg[7][23]  ( .D(n651), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][23] ) );
  DFFARX1 \regfile_reg[8][23]  ( .D(n650), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][23] ) );
  DFFARX1 \regfile_reg[9][23]  ( .D(n649), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][23] ) );
  DFFARX1 \regfile_reg[10][23]  ( .D(n648), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][23] ) );
  DFFARX1 \regfile_reg[11][23]  ( .D(n647), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][23] ) );
  DFFARX1 \regfile_reg[12][23]  ( .D(n646), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][23] ) );
  DFFARX1 \regfile_reg[13][23]  ( .D(n645), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][23] ) );
  DFFARX1 \regfile_reg[14][23]  ( .D(n644), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][23] ) );
  DFFARX1 \regfile_reg[15][23]  ( .D(n643), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][23] ) );
  DFFX1 \AluOut_reg[22]  ( .D(n642), .CLK(clk), .Q(AluOut[22]), .QN(n238) );
  DFFARX1 \regfile_reg[0][22]  ( .D(n641), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][22] ) );
  DFFARX1 \regfile_reg[1][22]  ( .D(n640), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][22] ) );
  DFFARX1 \regfile_reg[2][22]  ( .D(n639), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][22] ) );
  DFFARX1 \regfile_reg[3][22]  ( .D(n638), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][22] ) );
  DFFARX1 \regfile_reg[4][22]  ( .D(n637), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][22] ) );
  DFFARX1 \regfile_reg[5][22]  ( .D(n636), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][22] ) );
  DFFARX1 \regfile_reg[6][22]  ( .D(n635), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][22] ) );
  DFFARX1 \regfile_reg[7][22]  ( .D(n634), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][22] ) );
  DFFARX1 \regfile_reg[8][22]  ( .D(n633), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][22] ) );
  DFFARX1 \regfile_reg[9][22]  ( .D(n632), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][22] ) );
  DFFARX1 \regfile_reg[10][22]  ( .D(n631), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][22] ) );
  DFFARX1 \regfile_reg[11][22]  ( .D(n630), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][22] ) );
  DFFARX1 \regfile_reg[12][22]  ( .D(n629), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][22] ) );
  DFFARX1 \regfile_reg[13][22]  ( .D(n628), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][22] ) );
  DFFARX1 \regfile_reg[14][22]  ( .D(n627), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][22] ) );
  DFFARX1 \regfile_reg[15][22]  ( .D(n626), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][22] ) );
  DFFX1 \AluOut_reg[21]  ( .D(n625), .CLK(clk), .Q(AluOut[21]), .QN(n237) );
  DFFARX1 \regfile_reg[0][21]  ( .D(n624), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][21] ) );
  DFFARX1 \regfile_reg[1][21]  ( .D(n623), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][21] ) );
  DFFARX1 \regfile_reg[2][21]  ( .D(n622), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][21] ) );
  DFFARX1 \regfile_reg[3][21]  ( .D(n621), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][21] ) );
  DFFARX1 \regfile_reg[4][21]  ( .D(n620), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][21] ) );
  DFFARX1 \regfile_reg[5][21]  ( .D(n619), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][21] ) );
  DFFARX1 \regfile_reg[6][21]  ( .D(n618), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][21] ) );
  DFFARX1 \regfile_reg[7][21]  ( .D(n617), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][21] ) );
  DFFARX1 \regfile_reg[8][21]  ( .D(n616), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][21] ) );
  DFFARX1 \regfile_reg[9][21]  ( .D(n615), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][21] ) );
  DFFARX1 \regfile_reg[10][21]  ( .D(n614), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][21] ) );
  DFFARX1 \regfile_reg[11][21]  ( .D(n613), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][21] ) );
  DFFARX1 \regfile_reg[12][21]  ( .D(n612), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][21] ) );
  DFFARX1 \regfile_reg[13][21]  ( .D(n611), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][21] ) );
  DFFARX1 \regfile_reg[14][21]  ( .D(n610), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][21] ) );
  DFFARX1 \regfile_reg[15][21]  ( .D(n609), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][21] ) );
  DFFX1 \AluOut_reg[20]  ( .D(n608), .CLK(clk), .Q(AluOut[20]), .QN(n236) );
  DFFARX1 \regfile_reg[0][20]  ( .D(n607), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][20] ) );
  DFFARX1 \regfile_reg[1][20]  ( .D(n606), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][20] ) );
  DFFARX1 \regfile_reg[2][20]  ( .D(n605), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][20] ) );
  DFFARX1 \regfile_reg[3][20]  ( .D(n604), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][20] ) );
  DFFARX1 \regfile_reg[4][20]  ( .D(n603), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][20] ) );
  DFFARX1 \regfile_reg[5][20]  ( .D(n602), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][20] ) );
  DFFARX1 \regfile_reg[6][20]  ( .D(n601), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][20] ) );
  DFFARX1 \regfile_reg[7][20]  ( .D(n600), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][20] ) );
  DFFARX1 \regfile_reg[8][20]  ( .D(n599), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][20] ) );
  DFFARX1 \regfile_reg[9][20]  ( .D(n598), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][20] ) );
  DFFARX1 \regfile_reg[10][20]  ( .D(n597), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][20] ) );
  DFFARX1 \regfile_reg[11][20]  ( .D(n596), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][20] ) );
  DFFARX1 \regfile_reg[12][20]  ( .D(n595), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][20] ) );
  DFFARX1 \regfile_reg[13][20]  ( .D(n594), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][20] ) );
  DFFARX1 \regfile_reg[14][20]  ( .D(n593), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][20] ) );
  DFFARX1 \regfile_reg[15][20]  ( .D(n592), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][20] ) );
  DFFX1 \AluOut_reg[19]  ( .D(n591), .CLK(clk), .Q(AluOut[19]), .QN(n235) );
  DFFARX1 \regfile_reg[0][19]  ( .D(n590), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][19] ) );
  DFFARX1 \regfile_reg[1][19]  ( .D(n589), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][19] ) );
  DFFARX1 \regfile_reg[2][19]  ( .D(n588), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][19] ) );
  DFFARX1 \regfile_reg[3][19]  ( .D(n587), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][19] ) );
  DFFARX1 \regfile_reg[4][19]  ( .D(n586), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][19] ) );
  DFFARX1 \regfile_reg[5][19]  ( .D(n585), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][19] ) );
  DFFARX1 \regfile_reg[6][19]  ( .D(n584), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][19] ) );
  DFFARX1 \regfile_reg[7][19]  ( .D(n583), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][19] ) );
  DFFARX1 \regfile_reg[8][19]  ( .D(n582), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][19] ) );
  DFFARX1 \regfile_reg[9][19]  ( .D(n581), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][19] ) );
  DFFARX1 \regfile_reg[10][19]  ( .D(n580), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][19] ) );
  DFFARX1 \regfile_reg[11][19]  ( .D(n579), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][19] ) );
  DFFARX1 \regfile_reg[12][19]  ( .D(n578), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][19] ) );
  DFFARX1 \regfile_reg[13][19]  ( .D(n577), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][19] ) );
  DFFARX1 \regfile_reg[14][19]  ( .D(n576), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][19] ) );
  DFFARX1 \regfile_reg[15][19]  ( .D(n575), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][19] ) );
  DFFX1 \AluOut_reg[18]  ( .D(n574), .CLK(clk), .Q(AluOut[18]), .QN(n234) );
  DFFARX1 \regfile_reg[0][18]  ( .D(n573), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][18] ) );
  DFFARX1 \regfile_reg[1][18]  ( .D(n572), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][18] ) );
  DFFARX1 \regfile_reg[2][18]  ( .D(n571), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][18] ) );
  DFFARX1 \regfile_reg[3][18]  ( .D(n570), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][18] ) );
  DFFARX1 \regfile_reg[4][18]  ( .D(n569), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][18] ) );
  DFFARX1 \regfile_reg[5][18]  ( .D(n568), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][18] ) );
  DFFARX1 \regfile_reg[6][18]  ( .D(n567), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][18] ) );
  DFFARX1 \regfile_reg[7][18]  ( .D(n566), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][18] ) );
  DFFARX1 \regfile_reg[8][18]  ( .D(n565), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][18] ) );
  DFFARX1 \regfile_reg[9][18]  ( .D(n564), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][18] ) );
  DFFARX1 \regfile_reg[10][18]  ( .D(n563), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][18] ) );
  DFFARX1 \regfile_reg[11][18]  ( .D(n562), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][18] ) );
  DFFARX1 \regfile_reg[12][18]  ( .D(n561), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][18] ) );
  DFFARX1 \regfile_reg[13][18]  ( .D(n560), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][18] ) );
  DFFARX1 \regfile_reg[14][18]  ( .D(n559), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][18] ) );
  DFFARX1 \regfile_reg[15][18]  ( .D(n558), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][18] ) );
  DFFX1 \AluOut_reg[17]  ( .D(n557), .CLK(clk), .Q(AluOut[17]), .QN(n233) );
  DFFARX1 \regfile_reg[0][17]  ( .D(n556), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][17] ) );
  DFFARX1 \regfile_reg[1][17]  ( .D(n555), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][17] ) );
  DFFARX1 \regfile_reg[2][17]  ( .D(n554), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][17] ) );
  DFFARX1 \regfile_reg[3][17]  ( .D(n553), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][17] ) );
  DFFARX1 \regfile_reg[4][17]  ( .D(n552), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][17] ) );
  DFFARX1 \regfile_reg[5][17]  ( .D(n551), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][17] ) );
  DFFARX1 \regfile_reg[6][17]  ( .D(n550), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][17] ) );
  DFFARX1 \regfile_reg[7][17]  ( .D(n549), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][17] ) );
  DFFARX1 \regfile_reg[8][17]  ( .D(n548), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][17] ) );
  DFFARX1 \regfile_reg[9][17]  ( .D(n547), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][17] ) );
  DFFARX1 \regfile_reg[10][17]  ( .D(n546), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][17] ) );
  DFFARX1 \regfile_reg[11][17]  ( .D(n545), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][17] ) );
  DFFARX1 \regfile_reg[12][17]  ( .D(n544), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][17] ) );
  DFFARX1 \regfile_reg[13][17]  ( .D(n543), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][17] ) );
  DFFARX1 \regfile_reg[14][17]  ( .D(n542), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][17] ) );
  DFFARX1 \regfile_reg[15][17]  ( .D(n541), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][17] ) );
  DFFX1 \AluOut_reg[16]  ( .D(n540), .CLK(clk), .Q(AluOut[16]), .QN(n232) );
  DFFARX1 \regfile_reg[0][16]  ( .D(n539), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][16] ) );
  DFFARX1 \regfile_reg[1][16]  ( .D(n538), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][16] ) );
  DFFARX1 \regfile_reg[2][16]  ( .D(n537), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][16] ) );
  DFFARX1 \regfile_reg[3][16]  ( .D(n536), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][16] ) );
  DFFARX1 \regfile_reg[4][16]  ( .D(n535), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][16] ) );
  DFFARX1 \regfile_reg[5][16]  ( .D(n534), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][16] ) );
  DFFARX1 \regfile_reg[6][16]  ( .D(n533), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][16] ) );
  DFFARX1 \regfile_reg[7][16]  ( .D(n532), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][16] ) );
  DFFARX1 \regfile_reg[8][16]  ( .D(n531), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][16] ) );
  DFFARX1 \regfile_reg[9][16]  ( .D(n530), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][16] ) );
  DFFARX1 \regfile_reg[10][16]  ( .D(n529), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][16] ) );
  DFFARX1 \regfile_reg[11][16]  ( .D(n528), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][16] ) );
  DFFARX1 \regfile_reg[12][16]  ( .D(n527), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][16] ) );
  DFFARX1 \regfile_reg[13][16]  ( .D(n526), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][16] ) );
  DFFARX1 \regfile_reg[14][16]  ( .D(n525), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][16] ) );
  DFFARX1 \regfile_reg[15][16]  ( .D(n524), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][16] ) );
  DFFX1 \AluOut_reg[15]  ( .D(n523), .CLK(clk), .Q(AluOut[15]), .QN(n231) );
  DFFARX1 \regfile_reg[0][15]  ( .D(n522), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][15] ) );
  DFFARX1 \regfile_reg[1][15]  ( .D(n521), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][15] ) );
  DFFARX1 \regfile_reg[2][15]  ( .D(n520), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][15] ) );
  DFFARX1 \regfile_reg[3][15]  ( .D(n519), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][15] ) );
  DFFARX1 \regfile_reg[4][15]  ( .D(n518), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][15] ) );
  DFFARX1 \regfile_reg[5][15]  ( .D(n517), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][15] ) );
  DFFARX1 \regfile_reg[6][15]  ( .D(n516), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][15] ) );
  DFFARX1 \regfile_reg[7][15]  ( .D(n515), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][15] ) );
  DFFARX1 \regfile_reg[8][15]  ( .D(n514), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][15] ) );
  DFFARX1 \regfile_reg[9][15]  ( .D(n513), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][15] ) );
  DFFARX1 \regfile_reg[10][15]  ( .D(n512), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][15] ) );
  DFFARX1 \regfile_reg[11][15]  ( .D(n511), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][15] ) );
  DFFARX1 \regfile_reg[12][15]  ( .D(n510), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][15] ) );
  DFFARX1 \regfile_reg[13][15]  ( .D(n509), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][15] ) );
  DFFARX1 \regfile_reg[14][15]  ( .D(n508), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][15] ) );
  DFFARX1 \regfile_reg[15][15]  ( .D(n507), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][15] ) );
  DFFX1 \AluOut_reg[14]  ( .D(n506), .CLK(clk), .Q(AluOut[14]), .QN(n230) );
  DFFARX1 \regfile_reg[0][14]  ( .D(n505), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][14] ) );
  DFFARX1 \regfile_reg[1][14]  ( .D(n504), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][14] ) );
  DFFARX1 \regfile_reg[2][14]  ( .D(n503), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][14] ) );
  DFFARX1 \regfile_reg[3][14]  ( .D(n502), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][14] ) );
  DFFARX1 \regfile_reg[4][14]  ( .D(n501), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][14] ) );
  DFFARX1 \regfile_reg[5][14]  ( .D(n500), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][14] ) );
  DFFARX1 \regfile_reg[6][14]  ( .D(n499), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][14] ) );
  DFFARX1 \regfile_reg[7][14]  ( .D(n498), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][14] ) );
  DFFARX1 \regfile_reg[8][14]  ( .D(n497), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][14] ) );
  DFFARX1 \regfile_reg[9][14]  ( .D(n496), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][14] ) );
  DFFARX1 \regfile_reg[10][14]  ( .D(n495), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][14] ) );
  DFFARX1 \regfile_reg[11][14]  ( .D(n494), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][14] ) );
  DFFARX1 \regfile_reg[12][14]  ( .D(n493), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][14] ) );
  DFFARX1 \regfile_reg[13][14]  ( .D(n492), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][14] ) );
  DFFARX1 \regfile_reg[14][14]  ( .D(n491), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][14] ) );
  DFFARX1 \regfile_reg[15][14]  ( .D(n490), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][14] ) );
  DFFX1 \AluOut_reg[13]  ( .D(n489), .CLK(clk), .Q(AluOut[13]), .QN(n229) );
  DFFARX1 \regfile_reg[0][13]  ( .D(n488), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][13] ) );
  DFFARX1 \regfile_reg[1][13]  ( .D(n487), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][13] ) );
  DFFARX1 \regfile_reg[2][13]  ( .D(n486), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][13] ) );
  DFFARX1 \regfile_reg[3][13]  ( .D(n485), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][13] ) );
  DFFARX1 \regfile_reg[4][13]  ( .D(n484), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][13] ) );
  DFFARX1 \regfile_reg[5][13]  ( .D(n483), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][13] ) );
  DFFARX1 \regfile_reg[6][13]  ( .D(n482), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][13] ) );
  DFFARX1 \regfile_reg[7][13]  ( .D(n481), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][13] ) );
  DFFARX1 \regfile_reg[8][13]  ( .D(n480), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][13] ) );
  DFFARX1 \regfile_reg[9][13]  ( .D(n479), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][13] ) );
  DFFARX1 \regfile_reg[10][13]  ( .D(n478), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][13] ) );
  DFFARX1 \regfile_reg[11][13]  ( .D(n477), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][13] ) );
  DFFARX1 \regfile_reg[12][13]  ( .D(n476), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][13] ) );
  DFFARX1 \regfile_reg[13][13]  ( .D(n475), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][13] ) );
  DFFARX1 \regfile_reg[14][13]  ( .D(n474), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][13] ) );
  DFFARX1 \regfile_reg[15][13]  ( .D(n473), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][13] ) );
  DFFX1 \AluOut_reg[12]  ( .D(n472), .CLK(clk), .Q(AluOut[12]), .QN(n228) );
  DFFARX1 \regfile_reg[0][12]  ( .D(n471), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][12] ) );
  DFFARX1 \regfile_reg[1][12]  ( .D(n470), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][12] ) );
  DFFARX1 \regfile_reg[2][12]  ( .D(n469), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][12] ) );
  DFFARX1 \regfile_reg[3][12]  ( .D(n468), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][12] ) );
  DFFARX1 \regfile_reg[4][12]  ( .D(n467), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][12] ) );
  DFFARX1 \regfile_reg[5][12]  ( .D(n466), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][12] ) );
  DFFARX1 \regfile_reg[6][12]  ( .D(n465), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][12] ) );
  DFFARX1 \regfile_reg[7][12]  ( .D(n464), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][12] ) );
  DFFARX1 \regfile_reg[8][12]  ( .D(n463), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][12] ) );
  DFFARX1 \regfile_reg[9][12]  ( .D(n462), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][12] ) );
  DFFARX1 \regfile_reg[10][12]  ( .D(n461), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][12] ) );
  DFFARX1 \regfile_reg[11][12]  ( .D(n460), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][12] ) );
  DFFARX1 \regfile_reg[12][12]  ( .D(n459), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][12] ) );
  DFFARX1 \regfile_reg[13][12]  ( .D(n458), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][12] ) );
  DFFARX1 \regfile_reg[14][12]  ( .D(n457), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][12] ) );
  DFFARX1 \regfile_reg[15][12]  ( .D(n456), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][12] ) );
  DFFX1 \AluOut_reg[11]  ( .D(n455), .CLK(clk), .Q(AluOut[11]), .QN(n227) );
  DFFARX1 \regfile_reg[0][11]  ( .D(n454), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][11] ) );
  DFFARX1 \regfile_reg[1][11]  ( .D(n453), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][11] ) );
  DFFARX1 \regfile_reg[2][11]  ( .D(n452), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][11] ) );
  DFFARX1 \regfile_reg[3][11]  ( .D(n451), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][11] ) );
  DFFARX1 \regfile_reg[4][11]  ( .D(n450), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][11] ) );
  DFFARX1 \regfile_reg[5][11]  ( .D(n449), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][11] ) );
  DFFARX1 \regfile_reg[6][11]  ( .D(n448), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][11] ) );
  DFFARX1 \regfile_reg[7][11]  ( .D(n447), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][11] ) );
  DFFARX1 \regfile_reg[8][11]  ( .D(n446), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][11] ) );
  DFFARX1 \regfile_reg[9][11]  ( .D(n445), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][11] ) );
  DFFARX1 \regfile_reg[10][11]  ( .D(n444), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][11] ) );
  DFFARX1 \regfile_reg[11][11]  ( .D(n443), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][11] ) );
  DFFARX1 \regfile_reg[12][11]  ( .D(n442), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][11] ) );
  DFFARX1 \regfile_reg[13][11]  ( .D(n441), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][11] ) );
  DFFARX1 \regfile_reg[14][11]  ( .D(n440), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][11] ) );
  DFFARX1 \regfile_reg[15][11]  ( .D(n439), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][11] ) );
  DFFX1 \AluOut_reg[10]  ( .D(n438), .CLK(clk), .Q(AluOut[10]), .QN(n226) );
  DFFARX1 \regfile_reg[0][10]  ( .D(n437), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][10] ) );
  DFFARX1 \regfile_reg[1][10]  ( .D(n436), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][10] ) );
  DFFARX1 \regfile_reg[2][10]  ( .D(n435), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][10] ) );
  DFFARX1 \regfile_reg[3][10]  ( .D(n434), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][10] ) );
  DFFARX1 \regfile_reg[4][10]  ( .D(n433), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][10] ) );
  DFFARX1 \regfile_reg[5][10]  ( .D(n432), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][10] ) );
  DFFARX1 \regfile_reg[6][10]  ( .D(n431), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][10] ) );
  DFFARX1 \regfile_reg[7][10]  ( .D(n430), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][10] ) );
  DFFARX1 \regfile_reg[8][10]  ( .D(n429), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][10] ) );
  DFFARX1 \regfile_reg[9][10]  ( .D(n428), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][10] ) );
  DFFARX1 \regfile_reg[10][10]  ( .D(n427), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][10] ) );
  DFFARX1 \regfile_reg[11][10]  ( .D(n426), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][10] ) );
  DFFARX1 \regfile_reg[12][10]  ( .D(n425), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][10] ) );
  DFFARX1 \regfile_reg[13][10]  ( .D(n424), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][10] ) );
  DFFARX1 \regfile_reg[14][10]  ( .D(n423), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][10] ) );
  DFFARX1 \regfile_reg[15][10]  ( .D(n422), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][10] ) );
  DFFX1 \AluOut_reg[9]  ( .D(n421), .CLK(clk), .Q(AluOut[9]), .QN(n225) );
  DFFARX1 \regfile_reg[0][9]  ( .D(n420), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][9] ) );
  DFFARX1 \regfile_reg[1][9]  ( .D(n419), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][9] ) );
  DFFARX1 \regfile_reg[2][9]  ( .D(n418), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][9] ) );
  DFFARX1 \regfile_reg[3][9]  ( .D(n417), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][9] ) );
  DFFARX1 \regfile_reg[4][9]  ( .D(n416), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][9] ) );
  DFFARX1 \regfile_reg[5][9]  ( .D(n415), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][9] ) );
  DFFARX1 \regfile_reg[6][9]  ( .D(n414), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][9] ) );
  DFFARX1 \regfile_reg[7][9]  ( .D(n413), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][9] ) );
  DFFARX1 \regfile_reg[8][9]  ( .D(n412), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][9] ) );
  DFFARX1 \regfile_reg[9][9]  ( .D(n411), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][9] ) );
  DFFARX1 \regfile_reg[10][9]  ( .D(n410), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][9] ) );
  DFFARX1 \regfile_reg[11][9]  ( .D(n409), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][9] ) );
  DFFARX1 \regfile_reg[12][9]  ( .D(n408), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][9] ) );
  DFFARX1 \regfile_reg[13][9]  ( .D(n407), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][9] ) );
  DFFARX1 \regfile_reg[14][9]  ( .D(n406), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][9] ) );
  DFFARX1 \regfile_reg[15][9]  ( .D(n405), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][9] ) );
  DFFX1 \AluOut_reg[8]  ( .D(n404), .CLK(clk), .Q(AluOut[8]), .QN(n224) );
  DFFARX1 \regfile_reg[0][8]  ( .D(n403), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][8] ) );
  DFFARX1 \regfile_reg[1][8]  ( .D(n402), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][8] ) );
  DFFARX1 \regfile_reg[2][8]  ( .D(n401), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][8] ) );
  DFFARX1 \regfile_reg[3][8]  ( .D(n400), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][8] ) );
  DFFARX1 \regfile_reg[4][8]  ( .D(n399), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][8] ) );
  DFFARX1 \regfile_reg[5][8]  ( .D(n398), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][8] ) );
  DFFARX1 \regfile_reg[6][8]  ( .D(n397), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][8] ) );
  DFFARX1 \regfile_reg[7][8]  ( .D(n396), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][8] ) );
  DFFARX1 \regfile_reg[8][8]  ( .D(n395), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][8] ) );
  DFFARX1 \regfile_reg[9][8]  ( .D(n394), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][8] ) );
  DFFARX1 \regfile_reg[10][8]  ( .D(n393), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][8] ) );
  DFFARX1 \regfile_reg[11][8]  ( .D(n392), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][8] ) );
  DFFARX1 \regfile_reg[12][8]  ( .D(n391), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][8] ) );
  DFFARX1 \regfile_reg[13][8]  ( .D(n390), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][8] ) );
  DFFARX1 \regfile_reg[14][8]  ( .D(n389), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][8] ) );
  DFFARX1 \regfile_reg[15][8]  ( .D(n388), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][8] ) );
  DFFX1 \AluOut_reg[7]  ( .D(n387), .CLK(clk), .Q(AluOut[7]), .QN(n223) );
  DFFARX1 \regfile_reg[0][7]  ( .D(n386), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][7] ) );
  DFFARX1 \regfile_reg[1][7]  ( .D(n385), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][7] ) );
  DFFARX1 \regfile_reg[2][7]  ( .D(n384), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][7] ) );
  DFFARX1 \regfile_reg[3][7]  ( .D(n383), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][7] ) );
  DFFARX1 \regfile_reg[4][7]  ( .D(n382), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][7] ) );
  DFFARX1 \regfile_reg[5][7]  ( .D(n381), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][7] ) );
  DFFARX1 \regfile_reg[6][7]  ( .D(n380), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][7] ) );
  DFFARX1 \regfile_reg[7][7]  ( .D(n379), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][7] ) );
  DFFARX1 \regfile_reg[8][7]  ( .D(n378), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][7] ) );
  DFFARX1 \regfile_reg[9][7]  ( .D(n377), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][7] ) );
  DFFARX1 \regfile_reg[10][7]  ( .D(n376), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][7] ) );
  DFFARX1 \regfile_reg[11][7]  ( .D(n375), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][7] ) );
  DFFARX1 \regfile_reg[12][7]  ( .D(n374), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][7] ) );
  DFFARX1 \regfile_reg[13][7]  ( .D(n373), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][7] ) );
  DFFARX1 \regfile_reg[14][7]  ( .D(n372), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][7] ) );
  DFFARX1 \regfile_reg[15][7]  ( .D(n371), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][7] ) );
  DFFX1 \AluOut_reg[6]  ( .D(n370), .CLK(clk), .Q(AluOut[6]), .QN(n222) );
  DFFARX1 \regfile_reg[0][6]  ( .D(n369), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][6] ) );
  DFFARX1 \regfile_reg[1][6]  ( .D(n368), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][6] ) );
  DFFARX1 \regfile_reg[2][6]  ( .D(n367), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][6] ) );
  DFFARX1 \regfile_reg[3][6]  ( .D(n366), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][6] ) );
  DFFARX1 \regfile_reg[4][6]  ( .D(n365), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][6] ) );
  DFFARX1 \regfile_reg[5][6]  ( .D(n364), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][6] ) );
  DFFARX1 \regfile_reg[6][6]  ( .D(n363), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][6] ) );
  DFFARX1 \regfile_reg[7][6]  ( .D(n362), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][6] ) );
  DFFARX1 \regfile_reg[8][6]  ( .D(n361), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][6] ) );
  DFFARX1 \regfile_reg[9][6]  ( .D(n360), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][6] ) );
  DFFARX1 \regfile_reg[10][6]  ( .D(n359), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][6] ) );
  DFFARX1 \regfile_reg[11][6]  ( .D(n358), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][6] ) );
  DFFARX1 \regfile_reg[12][6]  ( .D(n357), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][6] ) );
  DFFARX1 \regfile_reg[13][6]  ( .D(n356), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][6] ) );
  DFFARX1 \regfile_reg[14][6]  ( .D(n355), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][6] ) );
  DFFARX1 \regfile_reg[15][6]  ( .D(n354), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][6] ) );
  DFFX1 \AluOut_reg[5]  ( .D(n353), .CLK(clk), .Q(AluOut[5]), .QN(n221) );
  DFFARX1 \regfile_reg[0][5]  ( .D(n352), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][5] ) );
  DFFARX1 \regfile_reg[1][5]  ( .D(n351), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][5] ) );
  DFFARX1 \regfile_reg[2][5]  ( .D(n350), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][5] ) );
  DFFARX1 \regfile_reg[3][5]  ( .D(n349), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][5] ) );
  DFFARX1 \regfile_reg[4][5]  ( .D(n348), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][5] ) );
  DFFARX1 \regfile_reg[5][5]  ( .D(n347), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][5] ) );
  DFFARX1 \regfile_reg[6][5]  ( .D(n346), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][5] ) );
  DFFARX1 \regfile_reg[7][5]  ( .D(n345), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][5] ) );
  DFFARX1 \regfile_reg[8][5]  ( .D(n344), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][5] ) );
  DFFARX1 \regfile_reg[9][5]  ( .D(n343), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][5] ) );
  DFFARX1 \regfile_reg[10][5]  ( .D(n342), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][5] ) );
  DFFARX1 \regfile_reg[11][5]  ( .D(n341), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][5] ) );
  DFFARX1 \regfile_reg[12][5]  ( .D(n340), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][5] ) );
  DFFARX1 \regfile_reg[13][5]  ( .D(n339), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][5] ) );
  DFFARX1 \regfile_reg[14][5]  ( .D(n338), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][5] ) );
  DFFARX1 \regfile_reg[15][5]  ( .D(n337), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][5] ) );
  DFFX1 \AluOut_reg[4]  ( .D(n336), .CLK(clk), .Q(AluOut[4]), .QN(n220) );
  DFFARX1 \regfile_reg[0][4]  ( .D(n335), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][4] ) );
  DFFARX1 \regfile_reg[1][4]  ( .D(n334), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][4] ) );
  DFFARX1 \regfile_reg[2][4]  ( .D(n333), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][4] ) );
  DFFARX1 \regfile_reg[3][4]  ( .D(n332), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][4] ) );
  DFFARX1 \regfile_reg[4][4]  ( .D(n331), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][4] ) );
  DFFARX1 \regfile_reg[5][4]  ( .D(n330), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][4] ) );
  DFFARX1 \regfile_reg[6][4]  ( .D(n329), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][4] ) );
  DFFARX1 \regfile_reg[7][4]  ( .D(n328), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][4] ) );
  DFFARX1 \regfile_reg[8][4]  ( .D(n327), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][4] ) );
  DFFARX1 \regfile_reg[9][4]  ( .D(n326), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][4] ) );
  DFFARX1 \regfile_reg[10][4]  ( .D(n325), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][4] ) );
  DFFARX1 \regfile_reg[11][4]  ( .D(n324), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][4] ) );
  DFFARX1 \regfile_reg[12][4]  ( .D(n323), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][4] ) );
  DFFARX1 \regfile_reg[13][4]  ( .D(n322), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][4] ) );
  DFFARX1 \regfile_reg[14][4]  ( .D(n321), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][4] ) );
  DFFASX1 \regfile_reg[15][4]  ( .D(n320), .CLK(clk), .SETB(rst), .Q(
        \regfile[15][4] ) );
  DFFX1 \AluOut_reg[3]  ( .D(n319), .CLK(clk), .Q(AluOut[3]), .QN(n219) );
  DFFARX1 \regfile_reg[0][3]  ( .D(n318), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][3] ) );
  DFFARX1 \regfile_reg[1][3]  ( .D(n317), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][3] ) );
  DFFARX1 \regfile_reg[2][3]  ( .D(n316), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][3] ) );
  DFFARX1 \regfile_reg[3][3]  ( .D(n315), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][3] ) );
  DFFARX1 \regfile_reg[4][3]  ( .D(n314), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][3] ) );
  DFFARX1 \regfile_reg[5][3]  ( .D(n313), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][3] ) );
  DFFARX1 \regfile_reg[6][3]  ( .D(n312), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][3] ) );
  DFFASX1 \regfile_reg[7][3]  ( .D(n311), .CLK(clk), .SETB(rst), .Q(
        \regfile[7][3] ) );
  DFFASX1 \regfile_reg[8][3]  ( .D(n310), .CLK(clk), .SETB(rst), .Q(
        \regfile[8][3] ) );
  DFFASX1 \regfile_reg[9][3]  ( .D(n309), .CLK(clk), .SETB(rst), .Q(
        \regfile[9][3] ) );
  DFFASX1 \regfile_reg[10][3]  ( .D(n308), .CLK(clk), .SETB(rst), .Q(
        \regfile[10][3] ) );
  DFFASX1 \regfile_reg[11][3]  ( .D(n307), .CLK(clk), .SETB(rst), .Q(
        \regfile[11][3] ) );
  DFFASX1 \regfile_reg[12][3]  ( .D(n306), .CLK(clk), .SETB(rst), .Q(
        \regfile[12][3] ) );
  DFFASX1 \regfile_reg[13][3]  ( .D(n305), .CLK(clk), .SETB(rst), .Q(
        \regfile[13][3] ) );
  DFFASX1 \regfile_reg[14][3]  ( .D(n304), .CLK(clk), .SETB(rst), .Q(
        \regfile[14][3] ) );
  DFFARX1 \regfile_reg[15][3]  ( .D(n303), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][3] ) );
  DFFX1 \AluOut_reg[2]  ( .D(n302), .CLK(clk), .Q(AluOut[2]), .QN(n218) );
  DFFARX1 \regfile_reg[0][2]  ( .D(n301), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][2] ) );
  DFFARX1 \regfile_reg[1][2]  ( .D(n300), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][2] ) );
  DFFARX1 \regfile_reg[2][2]  ( .D(n299), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][2] ) );
  DFFASX1 \regfile_reg[3][2]  ( .D(n298), .CLK(clk), .SETB(rst), .Q(
        \regfile[3][2] ) );
  DFFASX1 \regfile_reg[4][2]  ( .D(n297), .CLK(clk), .SETB(rst), .Q(
        \regfile[4][2] ) );
  DFFASX1 \regfile_reg[5][2]  ( .D(n296), .CLK(clk), .SETB(rst), .Q(
        \regfile[5][2] ) );
  DFFASX1 \regfile_reg[6][2]  ( .D(n295), .CLK(clk), .SETB(rst), .Q(
        \regfile[6][2] ) );
  DFFARX1 \regfile_reg[7][2]  ( .D(n294), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][2] ) );
  DFFARX1 \regfile_reg[8][2]  ( .D(n293), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][2] ) );
  DFFARX1 \regfile_reg[9][2]  ( .D(n292), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][2] ) );
  DFFARX1 \regfile_reg[10][2]  ( .D(n291), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][2] ) );
  DFFASX1 \regfile_reg[11][2]  ( .D(n290), .CLK(clk), .SETB(rst), .Q(
        \regfile[11][2] ) );
  DFFASX1 \regfile_reg[12][2]  ( .D(n289), .CLK(clk), .SETB(rst), .Q(
        \regfile[12][2] ) );
  DFFASX1 \regfile_reg[13][2]  ( .D(n288), .CLK(clk), .SETB(rst), .Q(
        \regfile[13][2] ) );
  DFFASX1 \regfile_reg[14][2]  ( .D(n287), .CLK(clk), .SETB(rst), .Q(
        \regfile[14][2] ) );
  DFFARX1 \regfile_reg[15][2]  ( .D(n286), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][2] ) );
  DFFX1 \AluOut_reg[1]  ( .D(n285), .CLK(clk), .Q(AluOut[1]), .QN(n217) );
  DFFARX1 \regfile_reg[0][1]  ( .D(n284), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][1] ) );
  DFFASX1 \regfile_reg[1][1]  ( .D(n283), .CLK(clk), .SETB(rst), .Q(
        \regfile[1][1] ) );
  DFFASX1 \regfile_reg[2][1]  ( .D(n282), .CLK(clk), .SETB(rst), .Q(
        \regfile[2][1] ) );
  DFFARX1 \regfile_reg[3][1]  ( .D(n281), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][1] ) );
  DFFARX1 \regfile_reg[4][1]  ( .D(n280), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][1] ) );
  DFFASX1 \regfile_reg[5][1]  ( .D(n279), .CLK(clk), .SETB(rst), .Q(
        \regfile[5][1] ) );
  DFFASX1 \regfile_reg[6][1]  ( .D(n278), .CLK(clk), .SETB(rst), .Q(
        \regfile[6][1] ) );
  DFFARX1 \regfile_reg[7][1]  ( .D(n277), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][1] ) );
  DFFARX1 \regfile_reg[8][1]  ( .D(n276), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][1] ) );
  DFFASX1 \regfile_reg[9][1]  ( .D(n275), .CLK(clk), .SETB(rst), .Q(
        \regfile[9][1] ) );
  DFFASX1 \regfile_reg[10][1]  ( .D(n274), .CLK(clk), .SETB(rst), .Q(
        \regfile[10][1] ) );
  DFFARX1 \regfile_reg[11][1]  ( .D(n273), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][1] ) );
  DFFARX1 \regfile_reg[12][1]  ( .D(n272), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][1] ) );
  DFFASX1 \regfile_reg[13][1]  ( .D(n271), .CLK(clk), .SETB(rst), .Q(
        \regfile[13][1] ) );
  DFFASX1 \regfile_reg[14][1]  ( .D(n270), .CLK(clk), .SETB(rst), .Q(
        \regfile[14][1] ) );
  DFFARX1 \regfile_reg[15][1]  ( .D(n269), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][1] ) );
  DFFX1 \AluOut_reg[0]  ( .D(n268), .CLK(clk), .Q(AluOut[0]), .QN(n216) );
  DFFASX1 \regfile_reg[0][0]  ( .D(n267), .CLK(clk), .SETB(rst), .Q(
        \regfile[0][0] ) );
  DFFARX1 \regfile_reg[1][0]  ( .D(n266), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][0] ) );
  DFFASX1 \regfile_reg[2][0]  ( .D(n265), .CLK(clk), .SETB(rst), .Q(
        \regfile[2][0] ) );
  DFFARX1 \regfile_reg[3][0]  ( .D(n264), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][0] ) );
  DFFASX1 \regfile_reg[4][0]  ( .D(n263), .CLK(clk), .SETB(rst), .Q(
        \regfile[4][0] ) );
  DFFARX1 \regfile_reg[5][0]  ( .D(n262), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][0] ) );
  DFFASX1 \regfile_reg[6][0]  ( .D(n261), .CLK(clk), .SETB(rst), .Q(
        \regfile[6][0] ) );
  DFFARX1 \regfile_reg[7][0]  ( .D(n260), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][0] ) );
  DFFASX1 \regfile_reg[8][0]  ( .D(n259), .CLK(clk), .SETB(rst), .Q(
        \regfile[8][0] ) );
  DFFARX1 \regfile_reg[9][0]  ( .D(n258), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][0] ) );
  DFFASX1 \regfile_reg[10][0]  ( .D(n257), .CLK(clk), .SETB(rst), .Q(
        \regfile[10][0] ) );
  DFFARX1 \regfile_reg[11][0]  ( .D(n256), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][0] ) );
  DFFASX1 \regfile_reg[12][0]  ( .D(n255), .CLK(clk), .SETB(rst), .Q(
        \regfile[12][0] ) );
  DFFARX1 \regfile_reg[13][0]  ( .D(n254), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][0] ) );
  DFFASX1 \regfile_reg[14][0]  ( .D(n253), .CLK(clk), .SETB(rst), .Q(
        \regfile[14][0] ) );
  DFFARX1 \regfile_reg[15][0]  ( .D(n252), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][0] ) );
  pipealu_DW01_addsub_0 r308 ( .A({1'b0, IFID_A}), .B({1'b0, IFID_B}), .CI(
        1'b0), .ADD_SUB(n1318), .SUM({N188, N187, N186, N185, N184, N183, N182, 
        N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, 
        N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, 
        N157, N156}) );
  OR2X1 U760 ( .IN1(n1285), .IN2(n1280), .Q(n798) );
  INVX0 U761 ( .INP(n798), .ZN(n801) );
  INVX0 U762 ( .INP(n798), .ZN(n802) );
  INVX0 U763 ( .INP(n798), .ZN(n803) );
  INVX0 U764 ( .INP(n798), .ZN(n804) );
  INVX2 U765 ( .INP(n1309), .ZN(n1318) );
  MUX41X1 U766 ( .IN1(\regfile[12][0] ), .IN3(\regfile[14][0] ), .IN2(
        \regfile[13][0] ), .IN4(\regfile[15][0] ), .S0(N16), .S1(N15), .Q(n805) );
  MUX41X1 U767 ( .IN1(\regfile[8][0] ), .IN3(\regfile[10][0] ), .IN2(
        \regfile[9][0] ), .IN4(\regfile[11][0] ), .S0(N16), .S1(N15), .Q(n806)
         );
  MUX41X1 U768 ( .IN1(\regfile[4][0] ), .IN3(\regfile[6][0] ), .IN2(
        \regfile[5][0] ), .IN4(\regfile[7][0] ), .S0(N16), .S1(N15), .Q(n807)
         );
  MUX41X1 U769 ( .IN1(\regfile[0][0] ), .IN3(\regfile[2][0] ), .IN2(
        \regfile[1][0] ), .IN4(\regfile[3][0] ), .S0(N16), .S1(N15), .Q(n808)
         );
  MUX41X1 U770 ( .IN1(n808), .IN3(n806), .IN2(n807), .IN4(n805), .S0(N18), 
        .S1(N17), .Q(IFID_A[0]) );
  MUX41X1 U771 ( .IN1(\regfile[12][1] ), .IN3(\regfile[14][1] ), .IN2(
        \regfile[13][1] ), .IN4(\regfile[15][1] ), .S0(N16), .S1(N15), .Q(n809) );
  MUX41X1 U772 ( .IN1(\regfile[8][1] ), .IN3(\regfile[10][1] ), .IN2(
        \regfile[9][1] ), .IN4(\regfile[11][1] ), .S0(N16), .S1(N15), .Q(n810)
         );
  MUX41X1 U773 ( .IN1(\regfile[4][1] ), .IN3(\regfile[6][1] ), .IN2(
        \regfile[5][1] ), .IN4(\regfile[7][1] ), .S0(N16), .S1(N15), .Q(n811)
         );
  MUX41X1 U774 ( .IN1(\regfile[0][1] ), .IN3(\regfile[2][1] ), .IN2(
        \regfile[1][1] ), .IN4(\regfile[3][1] ), .S0(N16), .S1(N15), .Q(n812)
         );
  MUX41X1 U775 ( .IN1(n812), .IN3(n810), .IN2(n811), .IN4(n809), .S0(N18), 
        .S1(N17), .Q(IFID_A[1]) );
  MUX41X1 U776 ( .IN1(\regfile[12][2] ), .IN3(\regfile[14][2] ), .IN2(
        \regfile[13][2] ), .IN4(\regfile[15][2] ), .S0(N16), .S1(N15), .Q(n813) );
  MUX41X1 U777 ( .IN1(\regfile[8][2] ), .IN3(\regfile[10][2] ), .IN2(
        \regfile[9][2] ), .IN4(\regfile[11][2] ), .S0(N16), .S1(N15), .Q(n814)
         );
  MUX41X1 U778 ( .IN1(\regfile[4][2] ), .IN3(\regfile[6][2] ), .IN2(
        \regfile[5][2] ), .IN4(\regfile[7][2] ), .S0(N16), .S1(N15), .Q(n815)
         );
  MUX41X1 U779 ( .IN1(\regfile[0][2] ), .IN3(\regfile[2][2] ), .IN2(
        \regfile[1][2] ), .IN4(\regfile[3][2] ), .S0(N16), .S1(N15), .Q(n816)
         );
  MUX41X1 U780 ( .IN1(n816), .IN3(n814), .IN2(n815), .IN4(n813), .S0(N18), 
        .S1(N17), .Q(IFID_A[2]) );
  MUX41X1 U781 ( .IN1(\regfile[12][3] ), .IN3(\regfile[14][3] ), .IN2(
        \regfile[13][3] ), .IN4(\regfile[15][3] ), .S0(N16), .S1(N15), .Q(n817) );
  MUX41X1 U782 ( .IN1(\regfile[8][3] ), .IN3(\regfile[10][3] ), .IN2(
        \regfile[9][3] ), .IN4(\regfile[11][3] ), .S0(N16), .S1(N15), .Q(n818)
         );
  MUX41X1 U783 ( .IN1(\regfile[4][3] ), .IN3(\regfile[6][3] ), .IN2(
        \regfile[5][3] ), .IN4(\regfile[7][3] ), .S0(N16), .S1(N15), .Q(n819)
         );
  MUX41X1 U784 ( .IN1(\regfile[0][3] ), .IN3(\regfile[2][3] ), .IN2(
        \regfile[1][3] ), .IN4(\regfile[3][3] ), .S0(N16), .S1(N15), .Q(n820)
         );
  MUX41X1 U785 ( .IN1(n820), .IN3(n818), .IN2(n819), .IN4(n817), .S0(N18), 
        .S1(N17), .Q(IFID_A[3]) );
  MUX41X1 U786 ( .IN1(\regfile[12][4] ), .IN3(\regfile[14][4] ), .IN2(
        \regfile[13][4] ), .IN4(\regfile[15][4] ), .S0(N16), .S1(N15), .Q(n821) );
  MUX41X1 U787 ( .IN1(\regfile[8][4] ), .IN3(\regfile[10][4] ), .IN2(
        \regfile[9][4] ), .IN4(\regfile[11][4] ), .S0(N16), .S1(N15), .Q(n822)
         );
  MUX41X1 U788 ( .IN1(\regfile[4][4] ), .IN3(\regfile[6][4] ), .IN2(
        \regfile[5][4] ), .IN4(\regfile[7][4] ), .S0(N16), .S1(N15), .Q(n823)
         );
  MUX41X1 U789 ( .IN1(\regfile[0][4] ), .IN3(\regfile[2][4] ), .IN2(
        \regfile[1][4] ), .IN4(\regfile[3][4] ), .S0(N16), .S1(N15), .Q(n824)
         );
  MUX41X1 U790 ( .IN1(n824), .IN3(n822), .IN2(n823), .IN4(n821), .S0(N18), 
        .S1(N17), .Q(IFID_A[4]) );
  MUX41X1 U791 ( .IN1(\regfile[12][5] ), .IN3(\regfile[14][5] ), .IN2(
        \regfile[13][5] ), .IN4(\regfile[15][5] ), .S0(N16), .S1(N15), .Q(n825) );
  MUX41X1 U792 ( .IN1(\regfile[8][5] ), .IN3(\regfile[10][5] ), .IN2(
        \regfile[9][5] ), .IN4(\regfile[11][5] ), .S0(N16), .S1(N15), .Q(n826)
         );
  MUX41X1 U793 ( .IN1(\regfile[4][5] ), .IN3(\regfile[6][5] ), .IN2(
        \regfile[5][5] ), .IN4(\regfile[7][5] ), .S0(N16), .S1(N15), .Q(n827)
         );
  MUX41X1 U794 ( .IN1(\regfile[0][5] ), .IN3(\regfile[2][5] ), .IN2(
        \regfile[1][5] ), .IN4(\regfile[3][5] ), .S0(N16), .S1(N15), .Q(n828)
         );
  MUX41X1 U795 ( .IN1(n828), .IN3(n826), .IN2(n827), .IN4(n825), .S0(N18), 
        .S1(N17), .Q(IFID_A[5]) );
  MUX41X1 U796 ( .IN1(\regfile[12][6] ), .IN3(\regfile[14][6] ), .IN2(
        \regfile[13][6] ), .IN4(\regfile[15][6] ), .S0(N16), .S1(N15), .Q(n829) );
  MUX41X1 U797 ( .IN1(\regfile[8][6] ), .IN3(\regfile[10][6] ), .IN2(
        \regfile[9][6] ), .IN4(\regfile[11][6] ), .S0(N16), .S1(N15), .Q(n830)
         );
  MUX41X1 U798 ( .IN1(\regfile[4][6] ), .IN3(\regfile[6][6] ), .IN2(
        \regfile[5][6] ), .IN4(\regfile[7][6] ), .S0(N16), .S1(N15), .Q(n831)
         );
  MUX41X1 U799 ( .IN1(\regfile[0][6] ), .IN3(\regfile[2][6] ), .IN2(
        \regfile[1][6] ), .IN4(\regfile[3][6] ), .S0(N16), .S1(N15), .Q(n832)
         );
  MUX41X1 U800 ( .IN1(n832), .IN3(n830), .IN2(n831), .IN4(n829), .S0(N18), 
        .S1(N17), .Q(IFID_A[6]) );
  MUX41X1 U801 ( .IN1(\regfile[12][7] ), .IN3(\regfile[14][7] ), .IN2(
        \regfile[13][7] ), .IN4(\regfile[15][7] ), .S0(N16), .S1(N15), .Q(n833) );
  MUX41X1 U802 ( .IN1(\regfile[8][7] ), .IN3(\regfile[10][7] ), .IN2(
        \regfile[9][7] ), .IN4(\regfile[11][7] ), .S0(N16), .S1(N15), .Q(n834)
         );
  MUX41X1 U803 ( .IN1(\regfile[4][7] ), .IN3(\regfile[6][7] ), .IN2(
        \regfile[5][7] ), .IN4(\regfile[7][7] ), .S0(N16), .S1(N15), .Q(n835)
         );
  MUX41X1 U804 ( .IN1(\regfile[0][7] ), .IN3(\regfile[2][7] ), .IN2(
        \regfile[1][7] ), .IN4(\regfile[3][7] ), .S0(N16), .S1(N15), .Q(n836)
         );
  MUX41X1 U805 ( .IN1(n836), .IN3(n834), .IN2(n835), .IN4(n833), .S0(N18), 
        .S1(N17), .Q(IFID_A[7]) );
  MUX41X1 U806 ( .IN1(\regfile[12][8] ), .IN3(\regfile[14][8] ), .IN2(
        \regfile[13][8] ), .IN4(\regfile[15][8] ), .S0(N16), .S1(N15), .Q(n837) );
  MUX41X1 U807 ( .IN1(\regfile[8][8] ), .IN3(\regfile[10][8] ), .IN2(
        \regfile[9][8] ), .IN4(\regfile[11][8] ), .S0(N16), .S1(N15), .Q(n838)
         );
  MUX41X1 U808 ( .IN1(\regfile[4][8] ), .IN3(\regfile[6][8] ), .IN2(
        \regfile[5][8] ), .IN4(\regfile[7][8] ), .S0(N16), .S1(N15), .Q(n839)
         );
  MUX41X1 U809 ( .IN1(\regfile[0][8] ), .IN3(\regfile[2][8] ), .IN2(
        \regfile[1][8] ), .IN4(\regfile[3][8] ), .S0(N16), .S1(N15), .Q(n840)
         );
  MUX41X1 U810 ( .IN1(n840), .IN3(n838), .IN2(n839), .IN4(n837), .S0(N18), 
        .S1(N17), .Q(IFID_A[8]) );
  MUX41X1 U811 ( .IN1(\regfile[12][9] ), .IN3(\regfile[14][9] ), .IN2(
        \regfile[13][9] ), .IN4(\regfile[15][9] ), .S0(N16), .S1(N15), .Q(n841) );
  MUX41X1 U812 ( .IN1(\regfile[8][9] ), .IN3(\regfile[10][9] ), .IN2(
        \regfile[9][9] ), .IN4(\regfile[11][9] ), .S0(N16), .S1(N15), .Q(n842)
         );
  MUX41X1 U813 ( .IN1(\regfile[4][9] ), .IN3(\regfile[6][9] ), .IN2(
        \regfile[5][9] ), .IN4(\regfile[7][9] ), .S0(N16), .S1(N15), .Q(n843)
         );
  MUX41X1 U814 ( .IN1(\regfile[0][9] ), .IN3(\regfile[2][9] ), .IN2(
        \regfile[1][9] ), .IN4(\regfile[3][9] ), .S0(N16), .S1(N15), .Q(n844)
         );
  MUX41X1 U815 ( .IN1(n844), .IN3(n842), .IN2(n843), .IN4(n841), .S0(N18), 
        .S1(N17), .Q(IFID_A[9]) );
  MUX41X1 U816 ( .IN1(\regfile[12][10] ), .IN3(\regfile[14][10] ), .IN2(
        \regfile[13][10] ), .IN4(\regfile[15][10] ), .S0(N16), .S1(N15), .Q(
        n845) );
  MUX41X1 U817 ( .IN1(\regfile[8][10] ), .IN3(\regfile[10][10] ), .IN2(
        \regfile[9][10] ), .IN4(\regfile[11][10] ), .S0(N16), .S1(N15), .Q(
        n846) );
  MUX41X1 U818 ( .IN1(\regfile[4][10] ), .IN3(\regfile[6][10] ), .IN2(
        \regfile[5][10] ), .IN4(\regfile[7][10] ), .S0(N16), .S1(N15), .Q(n847) );
  MUX41X1 U819 ( .IN1(\regfile[0][10] ), .IN3(\regfile[2][10] ), .IN2(
        \regfile[1][10] ), .IN4(\regfile[3][10] ), .S0(N16), .S1(N15), .Q(n848) );
  MUX41X1 U820 ( .IN1(n848), .IN3(n846), .IN2(n847), .IN4(n845), .S0(N18), 
        .S1(N17), .Q(IFID_A[10]) );
  MUX41X1 U821 ( .IN1(\regfile[12][11] ), .IN3(\regfile[14][11] ), .IN2(
        \regfile[13][11] ), .IN4(\regfile[15][11] ), .S0(N16), .S1(N15), .Q(
        n849) );
  MUX41X1 U822 ( .IN1(\regfile[8][11] ), .IN3(\regfile[10][11] ), .IN2(
        \regfile[9][11] ), .IN4(\regfile[11][11] ), .S0(N16), .S1(N15), .Q(
        n850) );
  MUX41X1 U823 ( .IN1(\regfile[4][11] ), .IN3(\regfile[6][11] ), .IN2(
        \regfile[5][11] ), .IN4(\regfile[7][11] ), .S0(N16), .S1(N15), .Q(n851) );
  MUX41X1 U824 ( .IN1(\regfile[0][11] ), .IN3(\regfile[2][11] ), .IN2(
        \regfile[1][11] ), .IN4(\regfile[3][11] ), .S0(N16), .S1(N15), .Q(n852) );
  MUX41X1 U825 ( .IN1(n852), .IN3(n850), .IN2(n851), .IN4(n849), .S0(N18), 
        .S1(N17), .Q(IFID_A[11]) );
  MUX41X1 U826 ( .IN1(\regfile[12][12] ), .IN3(\regfile[14][12] ), .IN2(
        \regfile[13][12] ), .IN4(\regfile[15][12] ), .S0(N16), .S1(N15), .Q(
        n853) );
  MUX41X1 U827 ( .IN1(\regfile[8][12] ), .IN3(\regfile[10][12] ), .IN2(
        \regfile[9][12] ), .IN4(\regfile[11][12] ), .S0(N16), .S1(N15), .Q(
        n854) );
  MUX41X1 U828 ( .IN1(\regfile[4][12] ), .IN3(\regfile[6][12] ), .IN2(
        \regfile[5][12] ), .IN4(\regfile[7][12] ), .S0(N16), .S1(N15), .Q(n855) );
  MUX41X1 U829 ( .IN1(\regfile[0][12] ), .IN3(\regfile[2][12] ), .IN2(
        \regfile[1][12] ), .IN4(\regfile[3][12] ), .S0(N16), .S1(N15), .Q(n856) );
  MUX41X1 U830 ( .IN1(n856), .IN3(n854), .IN2(n855), .IN4(n853), .S0(N18), 
        .S1(N17), .Q(IFID_A[12]) );
  MUX41X1 U831 ( .IN1(\regfile[12][13] ), .IN3(\regfile[14][13] ), .IN2(
        \regfile[13][13] ), .IN4(\regfile[15][13] ), .S0(N16), .S1(N15), .Q(
        n857) );
  MUX41X1 U832 ( .IN1(\regfile[8][13] ), .IN3(\regfile[10][13] ), .IN2(
        \regfile[9][13] ), .IN4(\regfile[11][13] ), .S0(N16), .S1(N15), .Q(
        n858) );
  MUX41X1 U833 ( .IN1(\regfile[4][13] ), .IN3(\regfile[6][13] ), .IN2(
        \regfile[5][13] ), .IN4(\regfile[7][13] ), .S0(N16), .S1(N15), .Q(n859) );
  MUX41X1 U834 ( .IN1(\regfile[0][13] ), .IN3(\regfile[2][13] ), .IN2(
        \regfile[1][13] ), .IN4(\regfile[3][13] ), .S0(N16), .S1(N15), .Q(n860) );
  MUX41X1 U835 ( .IN1(n860), .IN3(n858), .IN2(n859), .IN4(n857), .S0(N18), 
        .S1(N17), .Q(IFID_A[13]) );
  MUX41X1 U836 ( .IN1(\regfile[12][14] ), .IN3(\regfile[14][14] ), .IN2(
        \regfile[13][14] ), .IN4(\regfile[15][14] ), .S0(N16), .S1(N15), .Q(
        n861) );
  MUX41X1 U837 ( .IN1(\regfile[8][14] ), .IN3(\regfile[10][14] ), .IN2(
        \regfile[9][14] ), .IN4(\regfile[11][14] ), .S0(N16), .S1(N15), .Q(
        n862) );
  MUX41X1 U838 ( .IN1(\regfile[4][14] ), .IN3(\regfile[6][14] ), .IN2(
        \regfile[5][14] ), .IN4(\regfile[7][14] ), .S0(N16), .S1(N15), .Q(n863) );
  MUX41X1 U839 ( .IN1(\regfile[0][14] ), .IN3(\regfile[2][14] ), .IN2(
        \regfile[1][14] ), .IN4(\regfile[3][14] ), .S0(N16), .S1(N15), .Q(n864) );
  MUX41X1 U840 ( .IN1(n864), .IN3(n862), .IN2(n863), .IN4(n861), .S0(N18), 
        .S1(N17), .Q(IFID_A[14]) );
  MUX41X1 U841 ( .IN1(\regfile[12][15] ), .IN3(\regfile[14][15] ), .IN2(
        \regfile[13][15] ), .IN4(\regfile[15][15] ), .S0(N16), .S1(N15), .Q(
        n865) );
  MUX41X1 U842 ( .IN1(\regfile[8][15] ), .IN3(\regfile[10][15] ), .IN2(
        \regfile[9][15] ), .IN4(\regfile[11][15] ), .S0(N16), .S1(N15), .Q(
        n866) );
  MUX41X1 U843 ( .IN1(\regfile[4][15] ), .IN3(\regfile[6][15] ), .IN2(
        \regfile[5][15] ), .IN4(\regfile[7][15] ), .S0(N16), .S1(N15), .Q(n867) );
  MUX41X1 U844 ( .IN1(\regfile[0][15] ), .IN3(\regfile[2][15] ), .IN2(
        \regfile[1][15] ), .IN4(\regfile[3][15] ), .S0(N16), .S1(N15), .Q(n868) );
  MUX41X1 U845 ( .IN1(n868), .IN3(n866), .IN2(n867), .IN4(n865), .S0(N18), 
        .S1(N17), .Q(IFID_A[15]) );
  MUX41X1 U846 ( .IN1(\regfile[12][16] ), .IN3(\regfile[14][16] ), .IN2(
        \regfile[13][16] ), .IN4(\regfile[15][16] ), .S0(N16), .S1(N15), .Q(
        n869) );
  MUX41X1 U847 ( .IN1(\regfile[8][16] ), .IN3(\regfile[10][16] ), .IN2(
        \regfile[9][16] ), .IN4(\regfile[11][16] ), .S0(N16), .S1(N15), .Q(
        n870) );
  MUX41X1 U848 ( .IN1(\regfile[4][16] ), .IN3(\regfile[6][16] ), .IN2(
        \regfile[5][16] ), .IN4(\regfile[7][16] ), .S0(N16), .S1(N15), .Q(n871) );
  MUX41X1 U849 ( .IN1(\regfile[0][16] ), .IN3(\regfile[2][16] ), .IN2(
        \regfile[1][16] ), .IN4(\regfile[3][16] ), .S0(N16), .S1(N15), .Q(n872) );
  MUX41X1 U850 ( .IN1(n872), .IN3(n870), .IN2(n871), .IN4(n869), .S0(N18), 
        .S1(N17), .Q(IFID_A[16]) );
  MUX41X1 U851 ( .IN1(\regfile[12][17] ), .IN3(\regfile[14][17] ), .IN2(
        \regfile[13][17] ), .IN4(\regfile[15][17] ), .S0(N16), .S1(N15), .Q(
        n873) );
  MUX41X1 U852 ( .IN1(\regfile[8][17] ), .IN3(\regfile[10][17] ), .IN2(
        \regfile[9][17] ), .IN4(\regfile[11][17] ), .S0(N16), .S1(N15), .Q(
        n874) );
  MUX41X1 U853 ( .IN1(\regfile[4][17] ), .IN3(\regfile[6][17] ), .IN2(
        \regfile[5][17] ), .IN4(\regfile[7][17] ), .S0(N16), .S1(N15), .Q(n875) );
  MUX41X1 U854 ( .IN1(\regfile[0][17] ), .IN3(\regfile[2][17] ), .IN2(
        \regfile[1][17] ), .IN4(\regfile[3][17] ), .S0(N16), .S1(N15), .Q(n876) );
  MUX41X1 U855 ( .IN1(n876), .IN3(n874), .IN2(n875), .IN4(n873), .S0(N18), 
        .S1(N17), .Q(IFID_A[17]) );
  MUX41X1 U856 ( .IN1(\regfile[12][18] ), .IN3(\regfile[14][18] ), .IN2(
        \regfile[13][18] ), .IN4(\regfile[15][18] ), .S0(N16), .S1(N15), .Q(
        n877) );
  MUX41X1 U857 ( .IN1(\regfile[8][18] ), .IN3(\regfile[10][18] ), .IN2(
        \regfile[9][18] ), .IN4(\regfile[11][18] ), .S0(N16), .S1(N15), .Q(
        n878) );
  MUX41X1 U858 ( .IN1(\regfile[4][18] ), .IN3(\regfile[6][18] ), .IN2(
        \regfile[5][18] ), .IN4(\regfile[7][18] ), .S0(N16), .S1(N15), .Q(n879) );
  MUX41X1 U859 ( .IN1(\regfile[0][18] ), .IN3(\regfile[2][18] ), .IN2(
        \regfile[1][18] ), .IN4(\regfile[3][18] ), .S0(N16), .S1(N15), .Q(n880) );
  MUX41X1 U860 ( .IN1(n880), .IN3(n878), .IN2(n879), .IN4(n877), .S0(N18), 
        .S1(N17), .Q(IFID_A[18]) );
  MUX41X1 U861 ( .IN1(\regfile[12][19] ), .IN3(\regfile[14][19] ), .IN2(
        \regfile[13][19] ), .IN4(\regfile[15][19] ), .S0(N16), .S1(N15), .Q(
        n881) );
  MUX41X1 U862 ( .IN1(\regfile[8][19] ), .IN3(\regfile[10][19] ), .IN2(
        \regfile[9][19] ), .IN4(\regfile[11][19] ), .S0(N16), .S1(N15), .Q(
        n882) );
  MUX41X1 U863 ( .IN1(\regfile[4][19] ), .IN3(\regfile[6][19] ), .IN2(
        \regfile[5][19] ), .IN4(\regfile[7][19] ), .S0(N16), .S1(N15), .Q(n883) );
  MUX41X1 U864 ( .IN1(\regfile[0][19] ), .IN3(\regfile[2][19] ), .IN2(
        \regfile[1][19] ), .IN4(\regfile[3][19] ), .S0(N16), .S1(N15), .Q(n884) );
  MUX41X1 U865 ( .IN1(n884), .IN3(n882), .IN2(n883), .IN4(n881), .S0(N18), 
        .S1(N17), .Q(IFID_A[19]) );
  MUX41X1 U866 ( .IN1(\regfile[12][20] ), .IN3(\regfile[14][20] ), .IN2(
        \regfile[13][20] ), .IN4(\regfile[15][20] ), .S0(N16), .S1(N15), .Q(
        n885) );
  MUX41X1 U867 ( .IN1(\regfile[8][20] ), .IN3(\regfile[10][20] ), .IN2(
        \regfile[9][20] ), .IN4(\regfile[11][20] ), .S0(N16), .S1(N15), .Q(
        n886) );
  MUX41X1 U868 ( .IN1(\regfile[4][20] ), .IN3(\regfile[6][20] ), .IN2(
        \regfile[5][20] ), .IN4(\regfile[7][20] ), .S0(N16), .S1(N15), .Q(n887) );
  MUX41X1 U869 ( .IN1(\regfile[0][20] ), .IN3(\regfile[2][20] ), .IN2(
        \regfile[1][20] ), .IN4(\regfile[3][20] ), .S0(N16), .S1(N15), .Q(n888) );
  MUX41X1 U870 ( .IN1(n888), .IN3(n886), .IN2(n887), .IN4(n885), .S0(N18), 
        .S1(N17), .Q(IFID_A[20]) );
  MUX41X1 U871 ( .IN1(\regfile[12][21] ), .IN3(\regfile[14][21] ), .IN2(
        \regfile[13][21] ), .IN4(\regfile[15][21] ), .S0(N16), .S1(N15), .Q(
        n889) );
  MUX41X1 U872 ( .IN1(\regfile[8][21] ), .IN3(\regfile[10][21] ), .IN2(
        \regfile[9][21] ), .IN4(\regfile[11][21] ), .S0(N16), .S1(N15), .Q(
        n890) );
  MUX41X1 U873 ( .IN1(\regfile[4][21] ), .IN3(\regfile[6][21] ), .IN2(
        \regfile[5][21] ), .IN4(\regfile[7][21] ), .S0(N16), .S1(N15), .Q(n891) );
  MUX41X1 U874 ( .IN1(\regfile[0][21] ), .IN3(\regfile[2][21] ), .IN2(
        \regfile[1][21] ), .IN4(\regfile[3][21] ), .S0(N16), .S1(N15), .Q(n892) );
  MUX41X1 U875 ( .IN1(n892), .IN3(n890), .IN2(n891), .IN4(n889), .S0(N18), 
        .S1(N17), .Q(IFID_A[21]) );
  MUX41X1 U876 ( .IN1(\regfile[12][22] ), .IN3(\regfile[14][22] ), .IN2(
        \regfile[13][22] ), .IN4(\regfile[15][22] ), .S0(N16), .S1(N15), .Q(
        n893) );
  MUX41X1 U877 ( .IN1(\regfile[8][22] ), .IN3(\regfile[10][22] ), .IN2(
        \regfile[9][22] ), .IN4(\regfile[11][22] ), .S0(N16), .S1(N15), .Q(
        n894) );
  MUX41X1 U878 ( .IN1(\regfile[4][22] ), .IN3(\regfile[6][22] ), .IN2(
        \regfile[5][22] ), .IN4(\regfile[7][22] ), .S0(N16), .S1(N15), .Q(n895) );
  MUX41X1 U879 ( .IN1(\regfile[0][22] ), .IN3(\regfile[2][22] ), .IN2(
        \regfile[1][22] ), .IN4(\regfile[3][22] ), .S0(N16), .S1(N15), .Q(n896) );
  MUX41X1 U880 ( .IN1(n896), .IN3(n894), .IN2(n895), .IN4(n893), .S0(N18), 
        .S1(N17), .Q(IFID_A[22]) );
  MUX41X1 U881 ( .IN1(\regfile[12][23] ), .IN3(\regfile[14][23] ), .IN2(
        \regfile[13][23] ), .IN4(\regfile[15][23] ), .S0(N16), .S1(N15), .Q(
        n897) );
  MUX41X1 U882 ( .IN1(\regfile[8][23] ), .IN3(\regfile[10][23] ), .IN2(
        \regfile[9][23] ), .IN4(\regfile[11][23] ), .S0(N16), .S1(N15), .Q(
        n898) );
  MUX41X1 U883 ( .IN1(\regfile[4][23] ), .IN3(\regfile[6][23] ), .IN2(
        \regfile[5][23] ), .IN4(\regfile[7][23] ), .S0(N16), .S1(N15), .Q(n899) );
  MUX41X1 U884 ( .IN1(\regfile[0][23] ), .IN3(\regfile[2][23] ), .IN2(
        \regfile[1][23] ), .IN4(\regfile[3][23] ), .S0(N16), .S1(N15), .Q(n900) );
  MUX41X1 U885 ( .IN1(n900), .IN3(n898), .IN2(n899), .IN4(n897), .S0(N18), 
        .S1(N17), .Q(IFID_A[23]) );
  MUX41X1 U886 ( .IN1(\regfile[12][24] ), .IN3(\regfile[14][24] ), .IN2(
        \regfile[13][24] ), .IN4(\regfile[15][24] ), .S0(N16), .S1(N15), .Q(
        n901) );
  MUX41X1 U887 ( .IN1(\regfile[8][24] ), .IN3(\regfile[10][24] ), .IN2(
        \regfile[9][24] ), .IN4(\regfile[11][24] ), .S0(N16), .S1(N15), .Q(
        n902) );
  MUX41X1 U888 ( .IN1(\regfile[4][24] ), .IN3(\regfile[6][24] ), .IN2(
        \regfile[5][24] ), .IN4(\regfile[7][24] ), .S0(N16), .S1(N15), .Q(n903) );
  MUX41X1 U889 ( .IN1(\regfile[0][24] ), .IN3(\regfile[2][24] ), .IN2(
        \regfile[1][24] ), .IN4(\regfile[3][24] ), .S0(N16), .S1(N15), .Q(n904) );
  MUX41X1 U890 ( .IN1(n904), .IN3(n902), .IN2(n903), .IN4(n901), .S0(N18), 
        .S1(N17), .Q(IFID_A[24]) );
  MUX41X1 U891 ( .IN1(\regfile[12][25] ), .IN3(\regfile[14][25] ), .IN2(
        \regfile[13][25] ), .IN4(\regfile[15][25] ), .S0(N16), .S1(N15), .Q(
        n905) );
  MUX41X1 U892 ( .IN1(\regfile[8][25] ), .IN3(\regfile[10][25] ), .IN2(
        \regfile[9][25] ), .IN4(\regfile[11][25] ), .S0(N16), .S1(N15), .Q(
        n906) );
  MUX41X1 U893 ( .IN1(\regfile[4][25] ), .IN3(\regfile[6][25] ), .IN2(
        \regfile[5][25] ), .IN4(\regfile[7][25] ), .S0(N16), .S1(N15), .Q(n907) );
  MUX41X1 U894 ( .IN1(\regfile[0][25] ), .IN3(\regfile[2][25] ), .IN2(
        \regfile[1][25] ), .IN4(\regfile[3][25] ), .S0(N16), .S1(N15), .Q(n908) );
  MUX41X1 U895 ( .IN1(n908), .IN3(n906), .IN2(n907), .IN4(n905), .S0(N18), 
        .S1(N17), .Q(IFID_A[25]) );
  MUX41X1 U896 ( .IN1(\regfile[12][26] ), .IN3(\regfile[14][26] ), .IN2(
        \regfile[13][26] ), .IN4(\regfile[15][26] ), .S0(N16), .S1(N15), .Q(
        n909) );
  MUX41X1 U897 ( .IN1(\regfile[8][26] ), .IN3(\regfile[10][26] ), .IN2(
        \regfile[9][26] ), .IN4(\regfile[11][26] ), .S0(N16), .S1(N15), .Q(
        n910) );
  MUX41X1 U898 ( .IN1(\regfile[4][26] ), .IN3(\regfile[6][26] ), .IN2(
        \regfile[5][26] ), .IN4(\regfile[7][26] ), .S0(N16), .S1(N15), .Q(n911) );
  MUX41X1 U899 ( .IN1(\regfile[0][26] ), .IN3(\regfile[2][26] ), .IN2(
        \regfile[1][26] ), .IN4(\regfile[3][26] ), .S0(N16), .S1(N15), .Q(n912) );
  MUX41X1 U900 ( .IN1(n912), .IN3(n910), .IN2(n911), .IN4(n909), .S0(N18), 
        .S1(N17), .Q(IFID_A[26]) );
  MUX41X1 U901 ( .IN1(\regfile[12][27] ), .IN3(\regfile[14][27] ), .IN2(
        \regfile[13][27] ), .IN4(\regfile[15][27] ), .S0(N16), .S1(N15), .Q(
        n913) );
  MUX41X1 U902 ( .IN1(\regfile[8][27] ), .IN3(\regfile[10][27] ), .IN2(
        \regfile[9][27] ), .IN4(\regfile[11][27] ), .S0(N16), .S1(N15), .Q(
        n914) );
  MUX41X1 U903 ( .IN1(\regfile[4][27] ), .IN3(\regfile[6][27] ), .IN2(
        \regfile[5][27] ), .IN4(\regfile[7][27] ), .S0(N16), .S1(N15), .Q(n915) );
  MUX41X1 U904 ( .IN1(\regfile[0][27] ), .IN3(\regfile[2][27] ), .IN2(
        \regfile[1][27] ), .IN4(\regfile[3][27] ), .S0(N16), .S1(N15), .Q(n916) );
  MUX41X1 U905 ( .IN1(n916), .IN3(n914), .IN2(n915), .IN4(n913), .S0(N18), 
        .S1(N17), .Q(IFID_A[27]) );
  MUX41X1 U906 ( .IN1(\regfile[12][28] ), .IN3(\regfile[14][28] ), .IN2(
        \regfile[13][28] ), .IN4(\regfile[15][28] ), .S0(N16), .S1(N15), .Q(
        n917) );
  MUX41X1 U907 ( .IN1(\regfile[8][28] ), .IN3(\regfile[10][28] ), .IN2(
        \regfile[9][28] ), .IN4(\regfile[11][28] ), .S0(N16), .S1(N15), .Q(
        n918) );
  MUX41X1 U908 ( .IN1(\regfile[4][28] ), .IN3(\regfile[6][28] ), .IN2(
        \regfile[5][28] ), .IN4(\regfile[7][28] ), .S0(N16), .S1(N15), .Q(n919) );
  MUX41X1 U909 ( .IN1(\regfile[0][28] ), .IN3(\regfile[2][28] ), .IN2(
        \regfile[1][28] ), .IN4(\regfile[3][28] ), .S0(N16), .S1(N15), .Q(n920) );
  MUX41X1 U910 ( .IN1(n920), .IN3(n918), .IN2(n919), .IN4(n917), .S0(N18), 
        .S1(N17), .Q(IFID_A[28]) );
  MUX41X1 U911 ( .IN1(\regfile[12][29] ), .IN3(\regfile[14][29] ), .IN2(
        \regfile[13][29] ), .IN4(\regfile[15][29] ), .S0(N16), .S1(N15), .Q(
        n921) );
  MUX41X1 U912 ( .IN1(\regfile[8][29] ), .IN3(\regfile[10][29] ), .IN2(
        \regfile[9][29] ), .IN4(\regfile[11][29] ), .S0(N16), .S1(N15), .Q(
        n922) );
  MUX41X1 U913 ( .IN1(\regfile[4][29] ), .IN3(\regfile[6][29] ), .IN2(
        \regfile[5][29] ), .IN4(\regfile[7][29] ), .S0(N16), .S1(N15), .Q(n923) );
  MUX41X1 U914 ( .IN1(\regfile[0][29] ), .IN3(\regfile[2][29] ), .IN2(
        \regfile[1][29] ), .IN4(\regfile[3][29] ), .S0(N16), .S1(N15), .Q(n924) );
  MUX41X1 U915 ( .IN1(n924), .IN3(n922), .IN2(n923), .IN4(n921), .S0(N18), 
        .S1(N17), .Q(IFID_A[29]) );
  MUX41X1 U916 ( .IN1(\regfile[12][30] ), .IN3(\regfile[14][30] ), .IN2(
        \regfile[13][30] ), .IN4(\regfile[15][30] ), .S0(N16), .S1(N15), .Q(
        n925) );
  MUX41X1 U917 ( .IN1(\regfile[8][30] ), .IN3(\regfile[10][30] ), .IN2(
        \regfile[9][30] ), .IN4(\regfile[11][30] ), .S0(N16), .S1(N15), .Q(
        n926) );
  MUX41X1 U918 ( .IN1(\regfile[4][30] ), .IN3(\regfile[6][30] ), .IN2(
        \regfile[5][30] ), .IN4(\regfile[7][30] ), .S0(N16), .S1(N15), .Q(n927) );
  MUX41X1 U919 ( .IN1(\regfile[0][30] ), .IN3(\regfile[2][30] ), .IN2(
        \regfile[1][30] ), .IN4(\regfile[3][30] ), .S0(N16), .S1(N15), .Q(n928) );
  MUX41X1 U920 ( .IN1(n928), .IN3(n926), .IN2(n927), .IN4(n925), .S0(N18), 
        .S1(N17), .Q(IFID_A[30]) );
  MUX41X1 U921 ( .IN1(\regfile[12][31] ), .IN3(\regfile[14][31] ), .IN2(
        \regfile[13][31] ), .IN4(\regfile[15][31] ), .S0(N16), .S1(N15), .Q(
        n929) );
  MUX41X1 U922 ( .IN1(\regfile[8][31] ), .IN3(\regfile[10][31] ), .IN2(
        \regfile[9][31] ), .IN4(\regfile[11][31] ), .S0(N16), .S1(N15), .Q(
        n930) );
  MUX41X1 U923 ( .IN1(\regfile[4][31] ), .IN3(\regfile[6][31] ), .IN2(
        \regfile[5][31] ), .IN4(\regfile[7][31] ), .S0(N16), .S1(N15), .Q(n931) );
  MUX41X1 U924 ( .IN1(\regfile[0][31] ), .IN3(\regfile[2][31] ), .IN2(
        \regfile[1][31] ), .IN4(\regfile[3][31] ), .S0(N16), .S1(N15), .Q(n932) );
  MUX41X1 U925 ( .IN1(n932), .IN3(n930), .IN2(n931), .IN4(n929), .S0(N18), 
        .S1(N17), .Q(IFID_A[31]) );
  MUX41X1 U926 ( .IN1(\regfile[12][0] ), .IN3(\regfile[14][0] ), .IN2(
        \regfile[13][0] ), .IN4(\regfile[15][0] ), .S0(N20), .S1(N19), .Q(n933) );
  MUX41X1 U927 ( .IN1(\regfile[8][0] ), .IN3(\regfile[10][0] ), .IN2(
        \regfile[9][0] ), .IN4(\regfile[11][0] ), .S0(N20), .S1(N19), .Q(n934)
         );
  MUX41X1 U928 ( .IN1(\regfile[4][0] ), .IN3(\regfile[6][0] ), .IN2(
        \regfile[5][0] ), .IN4(\regfile[7][0] ), .S0(N20), .S1(N19), .Q(n935)
         );
  MUX41X1 U929 ( .IN1(\regfile[0][0] ), .IN3(\regfile[2][0] ), .IN2(
        \regfile[1][0] ), .IN4(\regfile[3][0] ), .S0(N20), .S1(N19), .Q(n936)
         );
  MUX41X1 U930 ( .IN1(n936), .IN3(n934), .IN2(n935), .IN4(n933), .S0(N22), 
        .S1(N21), .Q(IFID_B[0]) );
  MUX41X1 U931 ( .IN1(\regfile[12][1] ), .IN3(\regfile[14][1] ), .IN2(
        \regfile[13][1] ), .IN4(\regfile[15][1] ), .S0(N20), .S1(N19), .Q(n937) );
  MUX41X1 U932 ( .IN1(\regfile[8][1] ), .IN3(\regfile[10][1] ), .IN2(
        \regfile[9][1] ), .IN4(\regfile[11][1] ), .S0(N20), .S1(N19), .Q(n938)
         );
  MUX41X1 U933 ( .IN1(\regfile[4][1] ), .IN3(\regfile[6][1] ), .IN2(
        \regfile[5][1] ), .IN4(\regfile[7][1] ), .S0(N20), .S1(N19), .Q(n939)
         );
  MUX41X1 U934 ( .IN1(\regfile[0][1] ), .IN3(\regfile[2][1] ), .IN2(
        \regfile[1][1] ), .IN4(\regfile[3][1] ), .S0(N20), .S1(N19), .Q(n940)
         );
  MUX41X1 U935 ( .IN1(n940), .IN3(n938), .IN2(n939), .IN4(n937), .S0(N22), 
        .S1(N21), .Q(IFID_B[1]) );
  MUX41X1 U936 ( .IN1(\regfile[12][2] ), .IN3(\regfile[14][2] ), .IN2(
        \regfile[13][2] ), .IN4(\regfile[15][2] ), .S0(N20), .S1(N19), .Q(n941) );
  MUX41X1 U937 ( .IN1(\regfile[8][2] ), .IN3(\regfile[10][2] ), .IN2(
        \regfile[9][2] ), .IN4(\regfile[11][2] ), .S0(N20), .S1(N19), .Q(n942)
         );
  MUX41X1 U938 ( .IN1(\regfile[4][2] ), .IN3(\regfile[6][2] ), .IN2(
        \regfile[5][2] ), .IN4(\regfile[7][2] ), .S0(N20), .S1(N19), .Q(n943)
         );
  MUX41X1 U939 ( .IN1(\regfile[0][2] ), .IN3(\regfile[2][2] ), .IN2(
        \regfile[1][2] ), .IN4(\regfile[3][2] ), .S0(N20), .S1(N19), .Q(n944)
         );
  MUX41X1 U940 ( .IN1(n944), .IN3(n942), .IN2(n943), .IN4(n941), .S0(N22), 
        .S1(N21), .Q(IFID_B[2]) );
  MUX41X1 U941 ( .IN1(\regfile[12][3] ), .IN3(\regfile[14][3] ), .IN2(
        \regfile[13][3] ), .IN4(\regfile[15][3] ), .S0(N20), .S1(N19), .Q(n945) );
  MUX41X1 U942 ( .IN1(\regfile[8][3] ), .IN3(\regfile[10][3] ), .IN2(
        \regfile[9][3] ), .IN4(\regfile[11][3] ), .S0(N20), .S1(N19), .Q(n946)
         );
  MUX41X1 U943 ( .IN1(\regfile[4][3] ), .IN3(\regfile[6][3] ), .IN2(
        \regfile[5][3] ), .IN4(\regfile[7][3] ), .S0(N20), .S1(N19), .Q(n947)
         );
  MUX41X1 U944 ( .IN1(\regfile[0][3] ), .IN3(\regfile[2][3] ), .IN2(
        \regfile[1][3] ), .IN4(\regfile[3][3] ), .S0(N20), .S1(N19), .Q(n948)
         );
  MUX41X1 U945 ( .IN1(n948), .IN3(n946), .IN2(n947), .IN4(n945), .S0(N22), 
        .S1(N21), .Q(IFID_B[3]) );
  MUX41X1 U946 ( .IN1(\regfile[12][4] ), .IN3(\regfile[14][4] ), .IN2(
        \regfile[13][4] ), .IN4(\regfile[15][4] ), .S0(N20), .S1(N19), .Q(n949) );
  MUX41X1 U947 ( .IN1(\regfile[8][4] ), .IN3(\regfile[10][4] ), .IN2(
        \regfile[9][4] ), .IN4(\regfile[11][4] ), .S0(N20), .S1(N19), .Q(n950)
         );
  MUX41X1 U948 ( .IN1(\regfile[4][4] ), .IN3(\regfile[6][4] ), .IN2(
        \regfile[5][4] ), .IN4(\regfile[7][4] ), .S0(N20), .S1(N19), .Q(n951)
         );
  MUX41X1 U949 ( .IN1(\regfile[0][4] ), .IN3(\regfile[2][4] ), .IN2(
        \regfile[1][4] ), .IN4(\regfile[3][4] ), .S0(N20), .S1(N19), .Q(n952)
         );
  MUX41X1 U950 ( .IN1(n952), .IN3(n950), .IN2(n951), .IN4(n949), .S0(N22), 
        .S1(N21), .Q(IFID_B[4]) );
  MUX41X1 U951 ( .IN1(\regfile[12][5] ), .IN3(\regfile[14][5] ), .IN2(
        \regfile[13][5] ), .IN4(\regfile[15][5] ), .S0(N20), .S1(N19), .Q(n953) );
  MUX41X1 U952 ( .IN1(\regfile[8][5] ), .IN3(\regfile[10][5] ), .IN2(
        \regfile[9][5] ), .IN4(\regfile[11][5] ), .S0(N20), .S1(N19), .Q(n954)
         );
  MUX41X1 U953 ( .IN1(\regfile[4][5] ), .IN3(\regfile[6][5] ), .IN2(
        \regfile[5][5] ), .IN4(\regfile[7][5] ), .S0(N20), .S1(N19), .Q(n955)
         );
  MUX41X1 U954 ( .IN1(\regfile[0][5] ), .IN3(\regfile[2][5] ), .IN2(
        \regfile[1][5] ), .IN4(\regfile[3][5] ), .S0(N20), .S1(N19), .Q(n956)
         );
  MUX41X1 U955 ( .IN1(n956), .IN3(n954), .IN2(n955), .IN4(n953), .S0(N22), 
        .S1(N21), .Q(IFID_B[5]) );
  MUX41X1 U956 ( .IN1(\regfile[12][6] ), .IN3(\regfile[14][6] ), .IN2(
        \regfile[13][6] ), .IN4(\regfile[15][6] ), .S0(N20), .S1(N19), .Q(n957) );
  MUX41X1 U957 ( .IN1(\regfile[8][6] ), .IN3(\regfile[10][6] ), .IN2(
        \regfile[9][6] ), .IN4(\regfile[11][6] ), .S0(N20), .S1(N19), .Q(n958)
         );
  MUX41X1 U958 ( .IN1(\regfile[4][6] ), .IN3(\regfile[6][6] ), .IN2(
        \regfile[5][6] ), .IN4(\regfile[7][6] ), .S0(N20), .S1(N19), .Q(n959)
         );
  MUX41X1 U959 ( .IN1(\regfile[0][6] ), .IN3(\regfile[2][6] ), .IN2(
        \regfile[1][6] ), .IN4(\regfile[3][6] ), .S0(N20), .S1(N19), .Q(n960)
         );
  MUX41X1 U960 ( .IN1(n960), .IN3(n958), .IN2(n959), .IN4(n957), .S0(N22), 
        .S1(N21), .Q(IFID_B[6]) );
  MUX41X1 U961 ( .IN1(\regfile[12][7] ), .IN3(\regfile[14][7] ), .IN2(
        \regfile[13][7] ), .IN4(\regfile[15][7] ), .S0(N20), .S1(N19), .Q(n961) );
  MUX41X1 U962 ( .IN1(\regfile[8][7] ), .IN3(\regfile[10][7] ), .IN2(
        \regfile[9][7] ), .IN4(\regfile[11][7] ), .S0(N20), .S1(N19), .Q(n962)
         );
  MUX41X1 U963 ( .IN1(\regfile[4][7] ), .IN3(\regfile[6][7] ), .IN2(
        \regfile[5][7] ), .IN4(\regfile[7][7] ), .S0(N20), .S1(N19), .Q(n963)
         );
  MUX41X1 U964 ( .IN1(\regfile[0][7] ), .IN3(\regfile[2][7] ), .IN2(
        \regfile[1][7] ), .IN4(\regfile[3][7] ), .S0(N20), .S1(N19), .Q(n964)
         );
  MUX41X1 U965 ( .IN1(n964), .IN3(n962), .IN2(n963), .IN4(n961), .S0(N22), 
        .S1(N21), .Q(IFID_B[7]) );
  MUX41X1 U966 ( .IN1(\regfile[12][8] ), .IN3(\regfile[14][8] ), .IN2(
        \regfile[13][8] ), .IN4(\regfile[15][8] ), .S0(N20), .S1(N19), .Q(n965) );
  MUX41X1 U967 ( .IN1(\regfile[8][8] ), .IN3(\regfile[10][8] ), .IN2(
        \regfile[9][8] ), .IN4(\regfile[11][8] ), .S0(N20), .S1(N19), .Q(n966)
         );
  MUX41X1 U968 ( .IN1(\regfile[4][8] ), .IN3(\regfile[6][8] ), .IN2(
        \regfile[5][8] ), .IN4(\regfile[7][8] ), .S0(N20), .S1(N19), .Q(n967)
         );
  MUX41X1 U969 ( .IN1(\regfile[0][8] ), .IN3(\regfile[2][8] ), .IN2(
        \regfile[1][8] ), .IN4(\regfile[3][8] ), .S0(N20), .S1(N19), .Q(n968)
         );
  MUX41X1 U970 ( .IN1(n968), .IN3(n966), .IN2(n967), .IN4(n965), .S0(N22), 
        .S1(N21), .Q(IFID_B[8]) );
  MUX41X1 U971 ( .IN1(\regfile[12][9] ), .IN3(\regfile[14][9] ), .IN2(
        \regfile[13][9] ), .IN4(\regfile[15][9] ), .S0(N20), .S1(N19), .Q(n969) );
  MUX41X1 U972 ( .IN1(\regfile[8][9] ), .IN3(\regfile[10][9] ), .IN2(
        \regfile[9][9] ), .IN4(\regfile[11][9] ), .S0(N20), .S1(N19), .Q(n970)
         );
  MUX41X1 U973 ( .IN1(\regfile[4][9] ), .IN3(\regfile[6][9] ), .IN2(
        \regfile[5][9] ), .IN4(\regfile[7][9] ), .S0(N20), .S1(N19), .Q(n971)
         );
  MUX41X1 U974 ( .IN1(\regfile[0][9] ), .IN3(\regfile[2][9] ), .IN2(
        \regfile[1][9] ), .IN4(\regfile[3][9] ), .S0(N20), .S1(N19), .Q(n972)
         );
  MUX41X1 U975 ( .IN1(n972), .IN3(n970), .IN2(n971), .IN4(n969), .S0(N22), 
        .S1(N21), .Q(IFID_B[9]) );
  MUX41X1 U976 ( .IN1(\regfile[12][10] ), .IN3(\regfile[14][10] ), .IN2(
        \regfile[13][10] ), .IN4(\regfile[15][10] ), .S0(N20), .S1(N19), .Q(
        n973) );
  MUX41X1 U977 ( .IN1(\regfile[8][10] ), .IN3(\regfile[10][10] ), .IN2(
        \regfile[9][10] ), .IN4(\regfile[11][10] ), .S0(N20), .S1(N19), .Q(
        n974) );
  MUX41X1 U978 ( .IN1(\regfile[4][10] ), .IN3(\regfile[6][10] ), .IN2(
        \regfile[5][10] ), .IN4(\regfile[7][10] ), .S0(N20), .S1(N19), .Q(n975) );
  MUX41X1 U979 ( .IN1(\regfile[0][10] ), .IN3(\regfile[2][10] ), .IN2(
        \regfile[1][10] ), .IN4(\regfile[3][10] ), .S0(N20), .S1(N19), .Q(n976) );
  MUX41X1 U980 ( .IN1(n976), .IN3(n974), .IN2(n975), .IN4(n973), .S0(N22), 
        .S1(N21), .Q(IFID_B[10]) );
  MUX41X1 U981 ( .IN1(\regfile[12][11] ), .IN3(\regfile[14][11] ), .IN2(
        \regfile[13][11] ), .IN4(\regfile[15][11] ), .S0(N20), .S1(N19), .Q(
        n977) );
  MUX41X1 U982 ( .IN1(\regfile[8][11] ), .IN3(\regfile[10][11] ), .IN2(
        \regfile[9][11] ), .IN4(\regfile[11][11] ), .S0(N20), .S1(N19), .Q(
        n978) );
  MUX41X1 U983 ( .IN1(\regfile[4][11] ), .IN3(\regfile[6][11] ), .IN2(
        \regfile[5][11] ), .IN4(\regfile[7][11] ), .S0(N20), .S1(N19), .Q(n979) );
  MUX41X1 U984 ( .IN1(\regfile[0][11] ), .IN3(\regfile[2][11] ), .IN2(
        \regfile[1][11] ), .IN4(\regfile[3][11] ), .S0(N20), .S1(N19), .Q(n980) );
  MUX41X1 U985 ( .IN1(n980), .IN3(n978), .IN2(n979), .IN4(n977), .S0(N22), 
        .S1(N21), .Q(IFID_B[11]) );
  MUX41X1 U986 ( .IN1(\regfile[12][12] ), .IN3(\regfile[14][12] ), .IN2(
        \regfile[13][12] ), .IN4(\regfile[15][12] ), .S0(N20), .S1(N19), .Q(
        n981) );
  MUX41X1 U987 ( .IN1(\regfile[8][12] ), .IN3(\regfile[10][12] ), .IN2(
        \regfile[9][12] ), .IN4(\regfile[11][12] ), .S0(N20), .S1(N19), .Q(
        n982) );
  MUX41X1 U988 ( .IN1(\regfile[4][12] ), .IN3(\regfile[6][12] ), .IN2(
        \regfile[5][12] ), .IN4(\regfile[7][12] ), .S0(N20), .S1(N19), .Q(n983) );
  MUX41X1 U989 ( .IN1(\regfile[0][12] ), .IN3(\regfile[2][12] ), .IN2(
        \regfile[1][12] ), .IN4(\regfile[3][12] ), .S0(N20), .S1(N19), .Q(n984) );
  MUX41X1 U990 ( .IN1(n984), .IN3(n982), .IN2(n983), .IN4(n981), .S0(N22), 
        .S1(N21), .Q(IFID_B[12]) );
  MUX41X1 U991 ( .IN1(\regfile[12][13] ), .IN3(\regfile[14][13] ), .IN2(
        \regfile[13][13] ), .IN4(\regfile[15][13] ), .S0(N20), .S1(N19), .Q(
        n985) );
  MUX41X1 U992 ( .IN1(\regfile[8][13] ), .IN3(\regfile[10][13] ), .IN2(
        \regfile[9][13] ), .IN4(\regfile[11][13] ), .S0(N20), .S1(N19), .Q(
        n986) );
  MUX41X1 U993 ( .IN1(\regfile[4][13] ), .IN3(\regfile[6][13] ), .IN2(
        \regfile[5][13] ), .IN4(\regfile[7][13] ), .S0(N20), .S1(N19), .Q(n987) );
  MUX41X1 U994 ( .IN1(\regfile[0][13] ), .IN3(\regfile[2][13] ), .IN2(
        \regfile[1][13] ), .IN4(\regfile[3][13] ), .S0(N20), .S1(N19), .Q(n988) );
  MUX41X1 U995 ( .IN1(n988), .IN3(n986), .IN2(n987), .IN4(n985), .S0(N22), 
        .S1(N21), .Q(IFID_B[13]) );
  MUX41X1 U996 ( .IN1(\regfile[12][14] ), .IN3(\regfile[14][14] ), .IN2(
        \regfile[13][14] ), .IN4(\regfile[15][14] ), .S0(N20), .S1(N19), .Q(
        n989) );
  MUX41X1 U997 ( .IN1(\regfile[8][14] ), .IN3(\regfile[10][14] ), .IN2(
        \regfile[9][14] ), .IN4(\regfile[11][14] ), .S0(N20), .S1(N19), .Q(
        n990) );
  MUX41X1 U998 ( .IN1(\regfile[4][14] ), .IN3(\regfile[6][14] ), .IN2(
        \regfile[5][14] ), .IN4(\regfile[7][14] ), .S0(N20), .S1(N19), .Q(n991) );
  MUX41X1 U999 ( .IN1(\regfile[0][14] ), .IN3(\regfile[2][14] ), .IN2(
        \regfile[1][14] ), .IN4(\regfile[3][14] ), .S0(N20), .S1(N19), .Q(n992) );
  MUX41X1 U1000 ( .IN1(n992), .IN3(n990), .IN2(n991), .IN4(n989), .S0(N22), 
        .S1(N21), .Q(IFID_B[14]) );
  MUX41X1 U1001 ( .IN1(\regfile[12][15] ), .IN3(\regfile[14][15] ), .IN2(
        \regfile[13][15] ), .IN4(\regfile[15][15] ), .S0(N20), .S1(N19), .Q(
        n993) );
  MUX41X1 U1002 ( .IN1(\regfile[8][15] ), .IN3(\regfile[10][15] ), .IN2(
        \regfile[9][15] ), .IN4(\regfile[11][15] ), .S0(N20), .S1(N19), .Q(
        n994) );
  MUX41X1 U1003 ( .IN1(\regfile[4][15] ), .IN3(\regfile[6][15] ), .IN2(
        \regfile[5][15] ), .IN4(\regfile[7][15] ), .S0(N20), .S1(N19), .Q(n995) );
  MUX41X1 U1004 ( .IN1(\regfile[0][15] ), .IN3(\regfile[2][15] ), .IN2(
        \regfile[1][15] ), .IN4(\regfile[3][15] ), .S0(N20), .S1(N19), .Q(n996) );
  MUX41X1 U1005 ( .IN1(n996), .IN3(n994), .IN2(n995), .IN4(n993), .S0(N22), 
        .S1(N21), .Q(IFID_B[15]) );
  MUX41X1 U1006 ( .IN1(\regfile[12][16] ), .IN3(\regfile[14][16] ), .IN2(
        \regfile[13][16] ), .IN4(\regfile[15][16] ), .S0(N20), .S1(N19), .Q(
        n997) );
  MUX41X1 U1007 ( .IN1(\regfile[8][16] ), .IN3(\regfile[10][16] ), .IN2(
        \regfile[9][16] ), .IN4(\regfile[11][16] ), .S0(N20), .S1(N19), .Q(
        n998) );
  MUX41X1 U1008 ( .IN1(\regfile[4][16] ), .IN3(\regfile[6][16] ), .IN2(
        \regfile[5][16] ), .IN4(\regfile[7][16] ), .S0(N20), .S1(N19), .Q(n999) );
  MUX41X1 U1009 ( .IN1(\regfile[0][16] ), .IN3(\regfile[2][16] ), .IN2(
        \regfile[1][16] ), .IN4(\regfile[3][16] ), .S0(N20), .S1(N19), .Q(
        n1000) );
  MUX41X1 U1010 ( .IN1(n1000), .IN3(n998), .IN2(n999), .IN4(n997), .S0(N22), 
        .S1(N21), .Q(IFID_B[16]) );
  MUX41X1 U1011 ( .IN1(\regfile[12][17] ), .IN3(\regfile[14][17] ), .IN2(
        \regfile[13][17] ), .IN4(\regfile[15][17] ), .S0(N20), .S1(N19), .Q(
        n1001) );
  MUX41X1 U1012 ( .IN1(\regfile[8][17] ), .IN3(\regfile[10][17] ), .IN2(
        \regfile[9][17] ), .IN4(\regfile[11][17] ), .S0(N20), .S1(N19), .Q(
        n1002) );
  MUX41X1 U1013 ( .IN1(\regfile[4][17] ), .IN3(\regfile[6][17] ), .IN2(
        \regfile[5][17] ), .IN4(\regfile[7][17] ), .S0(N20), .S1(N19), .Q(
        n1003) );
  MUX41X1 U1014 ( .IN1(\regfile[0][17] ), .IN3(\regfile[2][17] ), .IN2(
        \regfile[1][17] ), .IN4(\regfile[3][17] ), .S0(N20), .S1(N19), .Q(
        n1004) );
  MUX41X1 U1015 ( .IN1(n1004), .IN3(n1002), .IN2(n1003), .IN4(n1001), .S0(N22), 
        .S1(N21), .Q(IFID_B[17]) );
  MUX41X1 U1016 ( .IN1(\regfile[12][18] ), .IN3(\regfile[14][18] ), .IN2(
        \regfile[13][18] ), .IN4(\regfile[15][18] ), .S0(N20), .S1(N19), .Q(
        n1005) );
  MUX41X1 U1017 ( .IN1(\regfile[8][18] ), .IN3(\regfile[10][18] ), .IN2(
        \regfile[9][18] ), .IN4(\regfile[11][18] ), .S0(N20), .S1(N19), .Q(
        n1006) );
  MUX41X1 U1018 ( .IN1(\regfile[4][18] ), .IN3(\regfile[6][18] ), .IN2(
        \regfile[5][18] ), .IN4(\regfile[7][18] ), .S0(N20), .S1(N19), .Q(
        n1007) );
  MUX41X1 U1019 ( .IN1(\regfile[0][18] ), .IN3(\regfile[2][18] ), .IN2(
        \regfile[1][18] ), .IN4(\regfile[3][18] ), .S0(N20), .S1(N19), .Q(
        n1008) );
  MUX41X1 U1020 ( .IN1(n1008), .IN3(n1006), .IN2(n1007), .IN4(n1005), .S0(N22), 
        .S1(N21), .Q(IFID_B[18]) );
  MUX41X1 U1021 ( .IN1(\regfile[12][19] ), .IN3(\regfile[14][19] ), .IN2(
        \regfile[13][19] ), .IN4(\regfile[15][19] ), .S0(N20), .S1(N19), .Q(
        n1009) );
  MUX41X1 U1022 ( .IN1(\regfile[8][19] ), .IN3(\regfile[10][19] ), .IN2(
        \regfile[9][19] ), .IN4(\regfile[11][19] ), .S0(N20), .S1(N19), .Q(
        n1010) );
  MUX41X1 U1023 ( .IN1(\regfile[4][19] ), .IN3(\regfile[6][19] ), .IN2(
        \regfile[5][19] ), .IN4(\regfile[7][19] ), .S0(N20), .S1(N19), .Q(
        n1011) );
  MUX41X1 U1024 ( .IN1(\regfile[0][19] ), .IN3(\regfile[2][19] ), .IN2(
        \regfile[1][19] ), .IN4(\regfile[3][19] ), .S0(N20), .S1(N19), .Q(
        n1012) );
  MUX41X1 U1025 ( .IN1(n1012), .IN3(n1010), .IN2(n1011), .IN4(n1009), .S0(N22), 
        .S1(N21), .Q(IFID_B[19]) );
  MUX41X1 U1026 ( .IN1(\regfile[12][20] ), .IN3(\regfile[14][20] ), .IN2(
        \regfile[13][20] ), .IN4(\regfile[15][20] ), .S0(N20), .S1(N19), .Q(
        n1013) );
  MUX41X1 U1027 ( .IN1(\regfile[8][20] ), .IN3(\regfile[10][20] ), .IN2(
        \regfile[9][20] ), .IN4(\regfile[11][20] ), .S0(N20), .S1(N19), .Q(
        n1014) );
  MUX41X1 U1028 ( .IN1(\regfile[4][20] ), .IN3(\regfile[6][20] ), .IN2(
        \regfile[5][20] ), .IN4(\regfile[7][20] ), .S0(N20), .S1(N19), .Q(
        n1015) );
  MUX41X1 U1029 ( .IN1(\regfile[0][20] ), .IN3(\regfile[2][20] ), .IN2(
        \regfile[1][20] ), .IN4(\regfile[3][20] ), .S0(N20), .S1(N19), .Q(
        n1016) );
  MUX41X1 U1030 ( .IN1(n1016), .IN3(n1014), .IN2(n1015), .IN4(n1013), .S0(N22), 
        .S1(N21), .Q(IFID_B[20]) );
  MUX41X1 U1031 ( .IN1(\regfile[12][21] ), .IN3(\regfile[14][21] ), .IN2(
        \regfile[13][21] ), .IN4(\regfile[15][21] ), .S0(N20), .S1(N19), .Q(
        n1017) );
  MUX41X1 U1032 ( .IN1(\regfile[8][21] ), .IN3(\regfile[10][21] ), .IN2(
        \regfile[9][21] ), .IN4(\regfile[11][21] ), .S0(N20), .S1(N19), .Q(
        n1018) );
  MUX41X1 U1033 ( .IN1(\regfile[4][21] ), .IN3(\regfile[6][21] ), .IN2(
        \regfile[5][21] ), .IN4(\regfile[7][21] ), .S0(N20), .S1(N19), .Q(
        n1019) );
  MUX41X1 U1034 ( .IN1(\regfile[0][21] ), .IN3(\regfile[2][21] ), .IN2(
        \regfile[1][21] ), .IN4(\regfile[3][21] ), .S0(N20), .S1(N19), .Q(
        n1020) );
  MUX41X1 U1035 ( .IN1(n1020), .IN3(n1018), .IN2(n1019), .IN4(n1017), .S0(N22), 
        .S1(N21), .Q(IFID_B[21]) );
  MUX41X1 U1036 ( .IN1(\regfile[12][22] ), .IN3(\regfile[14][22] ), .IN2(
        \regfile[13][22] ), .IN4(\regfile[15][22] ), .S0(N20), .S1(N19), .Q(
        n1021) );
  MUX41X1 U1037 ( .IN1(\regfile[8][22] ), .IN3(\regfile[10][22] ), .IN2(
        \regfile[9][22] ), .IN4(\regfile[11][22] ), .S0(N20), .S1(N19), .Q(
        n1022) );
  MUX41X1 U1038 ( .IN1(\regfile[4][22] ), .IN3(\regfile[6][22] ), .IN2(
        \regfile[5][22] ), .IN4(\regfile[7][22] ), .S0(N20), .S1(N19), .Q(
        n1023) );
  MUX41X1 U1039 ( .IN1(\regfile[0][22] ), .IN3(\regfile[2][22] ), .IN2(
        \regfile[1][22] ), .IN4(\regfile[3][22] ), .S0(N20), .S1(N19), .Q(
        n1024) );
  MUX41X1 U1040 ( .IN1(n1024), .IN3(n1022), .IN2(n1023), .IN4(n1021), .S0(N22), 
        .S1(N21), .Q(IFID_B[22]) );
  MUX41X1 U1041 ( .IN1(\regfile[12][23] ), .IN3(\regfile[14][23] ), .IN2(
        \regfile[13][23] ), .IN4(\regfile[15][23] ), .S0(N20), .S1(N19), .Q(
        n1025) );
  MUX41X1 U1042 ( .IN1(\regfile[8][23] ), .IN3(\regfile[10][23] ), .IN2(
        \regfile[9][23] ), .IN4(\regfile[11][23] ), .S0(N20), .S1(N19), .Q(
        n1026) );
  MUX41X1 U1043 ( .IN1(\regfile[4][23] ), .IN3(\regfile[6][23] ), .IN2(
        \regfile[5][23] ), .IN4(\regfile[7][23] ), .S0(N20), .S1(N19), .Q(
        n1027) );
  MUX41X1 U1044 ( .IN1(\regfile[0][23] ), .IN3(\regfile[2][23] ), .IN2(
        \regfile[1][23] ), .IN4(\regfile[3][23] ), .S0(N20), .S1(N19), .Q(
        n1028) );
  MUX41X1 U1045 ( .IN1(n1028), .IN3(n1026), .IN2(n1027), .IN4(n1025), .S0(N22), 
        .S1(N21), .Q(IFID_B[23]) );
  MUX41X1 U1046 ( .IN1(\regfile[12][24] ), .IN3(\regfile[14][24] ), .IN2(
        \regfile[13][24] ), .IN4(\regfile[15][24] ), .S0(N20), .S1(N19), .Q(
        n1029) );
  MUX41X1 U1047 ( .IN1(\regfile[8][24] ), .IN3(\regfile[10][24] ), .IN2(
        \regfile[9][24] ), .IN4(\regfile[11][24] ), .S0(N20), .S1(N19), .Q(
        n1030) );
  MUX41X1 U1048 ( .IN1(\regfile[4][24] ), .IN3(\regfile[6][24] ), .IN2(
        \regfile[5][24] ), .IN4(\regfile[7][24] ), .S0(N20), .S1(N19), .Q(
        n1031) );
  MUX41X1 U1049 ( .IN1(\regfile[0][24] ), .IN3(\regfile[2][24] ), .IN2(
        \regfile[1][24] ), .IN4(\regfile[3][24] ), .S0(N20), .S1(N19), .Q(
        n1032) );
  MUX41X1 U1050 ( .IN1(n1032), .IN3(n1030), .IN2(n1031), .IN4(n1029), .S0(N22), 
        .S1(N21), .Q(IFID_B[24]) );
  MUX41X1 U1051 ( .IN1(\regfile[12][25] ), .IN3(\regfile[14][25] ), .IN2(
        \regfile[13][25] ), .IN4(\regfile[15][25] ), .S0(N20), .S1(N19), .Q(
        n1033) );
  MUX41X1 U1052 ( .IN1(\regfile[8][25] ), .IN3(\regfile[10][25] ), .IN2(
        \regfile[9][25] ), .IN4(\regfile[11][25] ), .S0(N20), .S1(N19), .Q(
        n1034) );
  MUX41X1 U1053 ( .IN1(\regfile[4][25] ), .IN3(\regfile[6][25] ), .IN2(
        \regfile[5][25] ), .IN4(\regfile[7][25] ), .S0(N20), .S1(N19), .Q(
        n1035) );
  MUX41X1 U1054 ( .IN1(\regfile[0][25] ), .IN3(\regfile[2][25] ), .IN2(
        \regfile[1][25] ), .IN4(\regfile[3][25] ), .S0(N20), .S1(N19), .Q(
        n1036) );
  MUX41X1 U1055 ( .IN1(n1036), .IN3(n1034), .IN2(n1035), .IN4(n1033), .S0(N22), 
        .S1(N21), .Q(IFID_B[25]) );
  MUX41X1 U1056 ( .IN1(\regfile[12][26] ), .IN3(\regfile[14][26] ), .IN2(
        \regfile[13][26] ), .IN4(\regfile[15][26] ), .S0(N20), .S1(N19), .Q(
        n1037) );
  MUX41X1 U1057 ( .IN1(\regfile[8][26] ), .IN3(\regfile[10][26] ), .IN2(
        \regfile[9][26] ), .IN4(\regfile[11][26] ), .S0(N20), .S1(N19), .Q(
        n1038) );
  MUX41X1 U1058 ( .IN1(\regfile[4][26] ), .IN3(\regfile[6][26] ), .IN2(
        \regfile[5][26] ), .IN4(\regfile[7][26] ), .S0(N20), .S1(N19), .Q(
        n1039) );
  MUX41X1 U1059 ( .IN1(\regfile[0][26] ), .IN3(\regfile[2][26] ), .IN2(
        \regfile[1][26] ), .IN4(\regfile[3][26] ), .S0(N20), .S1(N19), .Q(
        n1040) );
  MUX41X1 U1060 ( .IN1(n1040), .IN3(n1038), .IN2(n1039), .IN4(n1037), .S0(N22), 
        .S1(N21), .Q(IFID_B[26]) );
  MUX41X1 U1061 ( .IN1(\regfile[12][27] ), .IN3(\regfile[14][27] ), .IN2(
        \regfile[13][27] ), .IN4(\regfile[15][27] ), .S0(N20), .S1(N19), .Q(
        n1041) );
  MUX41X1 U1062 ( .IN1(\regfile[8][27] ), .IN3(\regfile[10][27] ), .IN2(
        \regfile[9][27] ), .IN4(\regfile[11][27] ), .S0(N20), .S1(N19), .Q(
        n1042) );
  MUX41X1 U1063 ( .IN1(\regfile[4][27] ), .IN3(\regfile[6][27] ), .IN2(
        \regfile[5][27] ), .IN4(\regfile[7][27] ), .S0(N20), .S1(N19), .Q(
        n1043) );
  MUX41X1 U1064 ( .IN1(\regfile[0][27] ), .IN3(\regfile[2][27] ), .IN2(
        \regfile[1][27] ), .IN4(\regfile[3][27] ), .S0(N20), .S1(N19), .Q(
        n1044) );
  MUX41X1 U1065 ( .IN1(n1044), .IN3(n1042), .IN2(n1043), .IN4(n1041), .S0(N22), 
        .S1(N21), .Q(IFID_B[27]) );
  MUX41X1 U1066 ( .IN1(\regfile[12][28] ), .IN3(\regfile[14][28] ), .IN2(
        \regfile[13][28] ), .IN4(\regfile[15][28] ), .S0(N20), .S1(N19), .Q(
        n1045) );
  MUX41X1 U1067 ( .IN1(\regfile[8][28] ), .IN3(\regfile[10][28] ), .IN2(
        \regfile[9][28] ), .IN4(\regfile[11][28] ), .S0(N20), .S1(N19), .Q(
        n1046) );
  MUX41X1 U1068 ( .IN1(\regfile[4][28] ), .IN3(\regfile[6][28] ), .IN2(
        \regfile[5][28] ), .IN4(\regfile[7][28] ), .S0(N20), .S1(N19), .Q(
        n1047) );
  MUX41X1 U1069 ( .IN1(\regfile[0][28] ), .IN3(\regfile[2][28] ), .IN2(
        \regfile[1][28] ), .IN4(\regfile[3][28] ), .S0(N20), .S1(N19), .Q(
        n1048) );
  MUX41X1 U1070 ( .IN1(n1048), .IN3(n1046), .IN2(n1047), .IN4(n1045), .S0(N22), 
        .S1(N21), .Q(IFID_B[28]) );
  MUX41X1 U1071 ( .IN1(\regfile[12][29] ), .IN3(\regfile[14][29] ), .IN2(
        \regfile[13][29] ), .IN4(\regfile[15][29] ), .S0(N20), .S1(N19), .Q(
        n1049) );
  MUX41X1 U1072 ( .IN1(\regfile[8][29] ), .IN3(\regfile[10][29] ), .IN2(
        \regfile[9][29] ), .IN4(\regfile[11][29] ), .S0(N20), .S1(N19), .Q(
        n1050) );
  MUX41X1 U1073 ( .IN1(\regfile[4][29] ), .IN3(\regfile[6][29] ), .IN2(
        \regfile[5][29] ), .IN4(\regfile[7][29] ), .S0(N20), .S1(N19), .Q(
        n1051) );
  MUX41X1 U1074 ( .IN1(\regfile[0][29] ), .IN3(\regfile[2][29] ), .IN2(
        \regfile[1][29] ), .IN4(\regfile[3][29] ), .S0(N20), .S1(N19), .Q(
        n1052) );
  MUX41X1 U1075 ( .IN1(n1052), .IN3(n1050), .IN2(n1051), .IN4(n1049), .S0(N22), 
        .S1(N21), .Q(IFID_B[29]) );
  MUX41X1 U1076 ( .IN1(\regfile[12][30] ), .IN3(\regfile[14][30] ), .IN2(
        \regfile[13][30] ), .IN4(\regfile[15][30] ), .S0(N20), .S1(N19), .Q(
        n1053) );
  MUX41X1 U1077 ( .IN1(\regfile[8][30] ), .IN3(\regfile[10][30] ), .IN2(
        \regfile[9][30] ), .IN4(\regfile[11][30] ), .S0(N20), .S1(N19), .Q(
        n1054) );
  MUX41X1 U1078 ( .IN1(\regfile[4][30] ), .IN3(\regfile[6][30] ), .IN2(
        \regfile[5][30] ), .IN4(\regfile[7][30] ), .S0(N20), .S1(N19), .Q(
        n1055) );
  MUX41X1 U1079 ( .IN1(\regfile[0][30] ), .IN3(\regfile[2][30] ), .IN2(
        \regfile[1][30] ), .IN4(\regfile[3][30] ), .S0(N20), .S1(N19), .Q(
        n1056) );
  MUX41X1 U1080 ( .IN1(n1056), .IN3(n1054), .IN2(n1055), .IN4(n1053), .S0(N22), 
        .S1(N21), .Q(IFID_B[30]) );
  MUX41X1 U1081 ( .IN1(\regfile[12][31] ), .IN3(\regfile[14][31] ), .IN2(
        \regfile[13][31] ), .IN4(\regfile[15][31] ), .S0(N20), .S1(N19), .Q(
        n1057) );
  MUX41X1 U1082 ( .IN1(\regfile[8][31] ), .IN3(\regfile[10][31] ), .IN2(
        \regfile[9][31] ), .IN4(\regfile[11][31] ), .S0(N20), .S1(N19), .Q(
        n1058) );
  MUX41X1 U1083 ( .IN1(\regfile[4][31] ), .IN3(\regfile[6][31] ), .IN2(
        \regfile[5][31] ), .IN4(\regfile[7][31] ), .S0(N20), .S1(N19), .Q(
        n1059) );
  MUX41X1 U1084 ( .IN1(\regfile[0][31] ), .IN3(\regfile[2][31] ), .IN2(
        \regfile[1][31] ), .IN4(\regfile[3][31] ), .S0(N20), .S1(N19), .Q(
        n1060) );
  MUX41X1 U1085 ( .IN1(n1060), .IN3(n1058), .IN2(n1059), .IN4(n1057), .S0(N22), 
        .S1(N21), .Q(IFID_B[31]) );
  AO221X1 U1086 ( .IN1(n1061), .IN2(AluOut[31]), .IN3(N187), .IN4(n1062), 
        .IN5(n1063), .Q(n795) );
  AO21X1 U1087 ( .IN1(n801), .IN2(IFID_A[31]), .IN3(n1064), .Q(n1063) );
  MUX21X1 U1088 ( .IN1(n1065), .IN2(n1066), .S(IFID_B[31]), .Q(n1064) );
  AO21X1 U1089 ( .IN1(IFID_A[31]), .IN2(n1067), .IN3(n804), .Q(n1066) );
  NOR2X0 U1090 ( .IN1(IFID_A[31]), .IN2(n1068), .QN(n1065) );
  MUX21X1 U1091 ( .IN1(\regfile[0][31] ), .IN2(AluOut[31]), .S(n1069), .Q(n794) );
  MUX21X1 U1092 ( .IN1(\regfile[1][31] ), .IN2(AluOut[31]), .S(n1070), .Q(n793) );
  MUX21X1 U1093 ( .IN1(\regfile[2][31] ), .IN2(AluOut[31]), .S(n1071), .Q(n792) );
  MUX21X1 U1094 ( .IN1(\regfile[3][31] ), .IN2(AluOut[31]), .S(n1072), .Q(n791) );
  MUX21X1 U1095 ( .IN1(\regfile[4][31] ), .IN2(AluOut[31]), .S(n1073), .Q(n790) );
  MUX21X1 U1096 ( .IN1(\regfile[5][31] ), .IN2(AluOut[31]), .S(n1074), .Q(n789) );
  MUX21X1 U1097 ( .IN1(\regfile[6][31] ), .IN2(AluOut[31]), .S(n1075), .Q(n788) );
  MUX21X1 U1098 ( .IN1(\regfile[7][31] ), .IN2(AluOut[31]), .S(n1076), .Q(n787) );
  MUX21X1 U1099 ( .IN1(\regfile[8][31] ), .IN2(AluOut[31]), .S(n1077), .Q(n786) );
  MUX21X1 U1100 ( .IN1(\regfile[9][31] ), .IN2(AluOut[31]), .S(n1078), .Q(n785) );
  MUX21X1 U1101 ( .IN1(\regfile[10][31] ), .IN2(AluOut[31]), .S(n1079), .Q(
        n784) );
  MUX21X1 U1102 ( .IN1(\regfile[11][31] ), .IN2(AluOut[31]), .S(n1080), .Q(
        n783) );
  MUX21X1 U1103 ( .IN1(\regfile[12][31] ), .IN2(AluOut[31]), .S(n1081), .Q(
        n782) );
  MUX21X1 U1104 ( .IN1(\regfile[13][31] ), .IN2(AluOut[31]), .S(n1082), .Q(
        n781) );
  MUX21X1 U1105 ( .IN1(\regfile[14][31] ), .IN2(AluOut[31]), .S(n1083), .Q(
        n780) );
  MUX21X1 U1106 ( .IN1(\regfile[15][31] ), .IN2(AluOut[31]), .S(n1084), .Q(
        n779) );
  AO221X1 U1107 ( .IN1(n1061), .IN2(AluOut[30]), .IN3(N186), .IN4(n1062), 
        .IN5(n1085), .Q(n778) );
  AO21X1 U1108 ( .IN1(IFID_A[30]), .IN2(n803), .IN3(n1086), .Q(n1085) );
  MUX21X1 U1109 ( .IN1(n1087), .IN2(n1088), .S(IFID_B[30]), .Q(n1086) );
  AO21X1 U1110 ( .IN1(IFID_A[30]), .IN2(n1067), .IN3(n803), .Q(n1088) );
  NOR2X0 U1111 ( .IN1(IFID_A[30]), .IN2(n1068), .QN(n1087) );
  MUX21X1 U1112 ( .IN1(\regfile[0][30] ), .IN2(AluOut[30]), .S(n1069), .Q(n777) );
  MUX21X1 U1113 ( .IN1(\regfile[1][30] ), .IN2(AluOut[30]), .S(n1070), .Q(n776) );
  MUX21X1 U1114 ( .IN1(\regfile[2][30] ), .IN2(AluOut[30]), .S(n1071), .Q(n775) );
  MUX21X1 U1115 ( .IN1(\regfile[3][30] ), .IN2(AluOut[30]), .S(n1072), .Q(n774) );
  MUX21X1 U1116 ( .IN1(\regfile[4][30] ), .IN2(AluOut[30]), .S(n1073), .Q(n773) );
  MUX21X1 U1117 ( .IN1(\regfile[5][30] ), .IN2(AluOut[30]), .S(n1074), .Q(n772) );
  MUX21X1 U1118 ( .IN1(\regfile[6][30] ), .IN2(AluOut[30]), .S(n1075), .Q(n771) );
  MUX21X1 U1119 ( .IN1(\regfile[7][30] ), .IN2(AluOut[30]), .S(n1076), .Q(n770) );
  MUX21X1 U1120 ( .IN1(\regfile[8][30] ), .IN2(AluOut[30]), .S(n1077), .Q(n769) );
  MUX21X1 U1121 ( .IN1(\regfile[9][30] ), .IN2(AluOut[30]), .S(n1078), .Q(n768) );
  MUX21X1 U1122 ( .IN1(\regfile[10][30] ), .IN2(AluOut[30]), .S(n1079), .Q(
        n767) );
  MUX21X1 U1123 ( .IN1(\regfile[11][30] ), .IN2(AluOut[30]), .S(n1080), .Q(
        n766) );
  MUX21X1 U1124 ( .IN1(\regfile[12][30] ), .IN2(AluOut[30]), .S(n1081), .Q(
        n765) );
  MUX21X1 U1125 ( .IN1(\regfile[13][30] ), .IN2(AluOut[30]), .S(n1082), .Q(
        n764) );
  MUX21X1 U1126 ( .IN1(\regfile[14][30] ), .IN2(AluOut[30]), .S(n1083), .Q(
        n763) );
  MUX21X1 U1127 ( .IN1(\regfile[15][30] ), .IN2(AluOut[30]), .S(n1084), .Q(
        n762) );
  AO221X1 U1128 ( .IN1(n1061), .IN2(AluOut[29]), .IN3(N185), .IN4(n1062), 
        .IN5(n1089), .Q(n761) );
  AO21X1 U1129 ( .IN1(IFID_A[29]), .IN2(n802), .IN3(n1090), .Q(n1089) );
  MUX21X1 U1130 ( .IN1(n1091), .IN2(n1092), .S(IFID_B[29]), .Q(n1090) );
  AO21X1 U1131 ( .IN1(IFID_A[29]), .IN2(n1067), .IN3(n802), .Q(n1092) );
  NOR2X0 U1132 ( .IN1(IFID_A[29]), .IN2(n1068), .QN(n1091) );
  MUX21X1 U1133 ( .IN1(\regfile[0][29] ), .IN2(AluOut[29]), .S(n1069), .Q(n760) );
  MUX21X1 U1134 ( .IN1(\regfile[1][29] ), .IN2(AluOut[29]), .S(n1070), .Q(n759) );
  MUX21X1 U1135 ( .IN1(\regfile[2][29] ), .IN2(AluOut[29]), .S(n1071), .Q(n758) );
  MUX21X1 U1136 ( .IN1(\regfile[3][29] ), .IN2(AluOut[29]), .S(n1072), .Q(n757) );
  MUX21X1 U1137 ( .IN1(\regfile[4][29] ), .IN2(AluOut[29]), .S(n1073), .Q(n756) );
  MUX21X1 U1138 ( .IN1(\regfile[5][29] ), .IN2(AluOut[29]), .S(n1074), .Q(n755) );
  MUX21X1 U1139 ( .IN1(\regfile[6][29] ), .IN2(AluOut[29]), .S(n1075), .Q(n754) );
  MUX21X1 U1140 ( .IN1(\regfile[7][29] ), .IN2(AluOut[29]), .S(n1076), .Q(n753) );
  MUX21X1 U1141 ( .IN1(\regfile[8][29] ), .IN2(AluOut[29]), .S(n1077), .Q(n752) );
  MUX21X1 U1142 ( .IN1(\regfile[9][29] ), .IN2(AluOut[29]), .S(n1078), .Q(n751) );
  MUX21X1 U1143 ( .IN1(\regfile[10][29] ), .IN2(AluOut[29]), .S(n1079), .Q(
        n750) );
  MUX21X1 U1144 ( .IN1(\regfile[11][29] ), .IN2(AluOut[29]), .S(n1080), .Q(
        n749) );
  MUX21X1 U1145 ( .IN1(\regfile[12][29] ), .IN2(AluOut[29]), .S(n1081), .Q(
        n748) );
  MUX21X1 U1146 ( .IN1(\regfile[13][29] ), .IN2(AluOut[29]), .S(n1082), .Q(
        n747) );
  MUX21X1 U1147 ( .IN1(\regfile[14][29] ), .IN2(AluOut[29]), .S(n1083), .Q(
        n746) );
  MUX21X1 U1148 ( .IN1(\regfile[15][29] ), .IN2(AluOut[29]), .S(n1084), .Q(
        n745) );
  AO221X1 U1149 ( .IN1(n1061), .IN2(AluOut[28]), .IN3(N184), .IN4(n1062), 
        .IN5(n1093), .Q(n744) );
  AO21X1 U1150 ( .IN1(IFID_A[28]), .IN2(n801), .IN3(n1094), .Q(n1093) );
  MUX21X1 U1151 ( .IN1(n1095), .IN2(n1096), .S(IFID_B[28]), .Q(n1094) );
  AO21X1 U1152 ( .IN1(IFID_A[28]), .IN2(n1067), .IN3(n801), .Q(n1096) );
  NOR2X0 U1153 ( .IN1(IFID_A[28]), .IN2(n1068), .QN(n1095) );
  MUX21X1 U1154 ( .IN1(\regfile[0][28] ), .IN2(AluOut[28]), .S(n1069), .Q(n743) );
  MUX21X1 U1155 ( .IN1(\regfile[1][28] ), .IN2(AluOut[28]), .S(n1070), .Q(n742) );
  MUX21X1 U1156 ( .IN1(\regfile[2][28] ), .IN2(AluOut[28]), .S(n1071), .Q(n741) );
  MUX21X1 U1157 ( .IN1(\regfile[3][28] ), .IN2(AluOut[28]), .S(n1072), .Q(n740) );
  MUX21X1 U1158 ( .IN1(\regfile[4][28] ), .IN2(AluOut[28]), .S(n1073), .Q(n739) );
  MUX21X1 U1159 ( .IN1(\regfile[5][28] ), .IN2(AluOut[28]), .S(n1074), .Q(n738) );
  MUX21X1 U1160 ( .IN1(\regfile[6][28] ), .IN2(AluOut[28]), .S(n1075), .Q(n737) );
  MUX21X1 U1161 ( .IN1(\regfile[7][28] ), .IN2(AluOut[28]), .S(n1076), .Q(n736) );
  MUX21X1 U1162 ( .IN1(\regfile[8][28] ), .IN2(AluOut[28]), .S(n1077), .Q(n735) );
  MUX21X1 U1163 ( .IN1(\regfile[9][28] ), .IN2(AluOut[28]), .S(n1078), .Q(n734) );
  MUX21X1 U1164 ( .IN1(\regfile[10][28] ), .IN2(AluOut[28]), .S(n1079), .Q(
        n733) );
  MUX21X1 U1165 ( .IN1(\regfile[11][28] ), .IN2(AluOut[28]), .S(n1080), .Q(
        n732) );
  MUX21X1 U1166 ( .IN1(\regfile[12][28] ), .IN2(AluOut[28]), .S(n1081), .Q(
        n731) );
  MUX21X1 U1167 ( .IN1(\regfile[13][28] ), .IN2(AluOut[28]), .S(n1082), .Q(
        n730) );
  MUX21X1 U1168 ( .IN1(\regfile[14][28] ), .IN2(AluOut[28]), .S(n1083), .Q(
        n729) );
  MUX21X1 U1169 ( .IN1(\regfile[15][28] ), .IN2(AluOut[28]), .S(n1084), .Q(
        n728) );
  AO221X1 U1170 ( .IN1(n1061), .IN2(AluOut[27]), .IN3(N183), .IN4(n1062), 
        .IN5(n1097), .Q(n727) );
  AO21X1 U1171 ( .IN1(IFID_A[27]), .IN2(n804), .IN3(n1098), .Q(n1097) );
  MUX21X1 U1172 ( .IN1(n1099), .IN2(n1100), .S(IFID_B[27]), .Q(n1098) );
  AO21X1 U1173 ( .IN1(IFID_A[27]), .IN2(n1067), .IN3(n804), .Q(n1100) );
  NOR2X0 U1174 ( .IN1(IFID_A[27]), .IN2(n1068), .QN(n1099) );
  MUX21X1 U1175 ( .IN1(\regfile[0][27] ), .IN2(AluOut[27]), .S(n1069), .Q(n726) );
  MUX21X1 U1176 ( .IN1(\regfile[1][27] ), .IN2(AluOut[27]), .S(n1070), .Q(n725) );
  MUX21X1 U1177 ( .IN1(\regfile[2][27] ), .IN2(AluOut[27]), .S(n1071), .Q(n724) );
  MUX21X1 U1178 ( .IN1(\regfile[3][27] ), .IN2(AluOut[27]), .S(n1072), .Q(n723) );
  MUX21X1 U1179 ( .IN1(\regfile[4][27] ), .IN2(AluOut[27]), .S(n1073), .Q(n722) );
  MUX21X1 U1180 ( .IN1(\regfile[5][27] ), .IN2(AluOut[27]), .S(n1074), .Q(n721) );
  MUX21X1 U1181 ( .IN1(\regfile[6][27] ), .IN2(AluOut[27]), .S(n1075), .Q(n720) );
  MUX21X1 U1182 ( .IN1(\regfile[7][27] ), .IN2(AluOut[27]), .S(n1076), .Q(n719) );
  MUX21X1 U1183 ( .IN1(\regfile[8][27] ), .IN2(AluOut[27]), .S(n1077), .Q(n718) );
  MUX21X1 U1184 ( .IN1(\regfile[9][27] ), .IN2(AluOut[27]), .S(n1078), .Q(n717) );
  MUX21X1 U1185 ( .IN1(\regfile[10][27] ), .IN2(AluOut[27]), .S(n1079), .Q(
        n716) );
  MUX21X1 U1186 ( .IN1(\regfile[11][27] ), .IN2(AluOut[27]), .S(n1080), .Q(
        n715) );
  MUX21X1 U1187 ( .IN1(\regfile[12][27] ), .IN2(AluOut[27]), .S(n1081), .Q(
        n714) );
  MUX21X1 U1188 ( .IN1(\regfile[13][27] ), .IN2(AluOut[27]), .S(n1082), .Q(
        n713) );
  MUX21X1 U1189 ( .IN1(\regfile[14][27] ), .IN2(AluOut[27]), .S(n1083), .Q(
        n712) );
  MUX21X1 U1190 ( .IN1(\regfile[15][27] ), .IN2(AluOut[27]), .S(n1084), .Q(
        n711) );
  AO221X1 U1191 ( .IN1(n1061), .IN2(AluOut[26]), .IN3(N182), .IN4(n1062), 
        .IN5(n1101), .Q(n710) );
  AO21X1 U1192 ( .IN1(IFID_A[26]), .IN2(n803), .IN3(n1102), .Q(n1101) );
  MUX21X1 U1193 ( .IN1(n1103), .IN2(n1104), .S(IFID_B[26]), .Q(n1102) );
  AO21X1 U1194 ( .IN1(IFID_A[26]), .IN2(n1067), .IN3(n803), .Q(n1104) );
  NOR2X0 U1195 ( .IN1(IFID_A[26]), .IN2(n1068), .QN(n1103) );
  MUX21X1 U1196 ( .IN1(\regfile[0][26] ), .IN2(AluOut[26]), .S(n1069), .Q(n709) );
  MUX21X1 U1197 ( .IN1(\regfile[1][26] ), .IN2(AluOut[26]), .S(n1070), .Q(n708) );
  MUX21X1 U1198 ( .IN1(\regfile[2][26] ), .IN2(AluOut[26]), .S(n1071), .Q(n707) );
  MUX21X1 U1199 ( .IN1(\regfile[3][26] ), .IN2(AluOut[26]), .S(n1072), .Q(n706) );
  MUX21X1 U1200 ( .IN1(\regfile[4][26] ), .IN2(AluOut[26]), .S(n1073), .Q(n705) );
  MUX21X1 U1201 ( .IN1(\regfile[5][26] ), .IN2(AluOut[26]), .S(n1074), .Q(n704) );
  MUX21X1 U1202 ( .IN1(\regfile[6][26] ), .IN2(AluOut[26]), .S(n1075), .Q(n703) );
  MUX21X1 U1203 ( .IN1(\regfile[7][26] ), .IN2(AluOut[26]), .S(n1076), .Q(n702) );
  MUX21X1 U1204 ( .IN1(\regfile[8][26] ), .IN2(AluOut[26]), .S(n1077), .Q(n701) );
  MUX21X1 U1205 ( .IN1(\regfile[9][26] ), .IN2(AluOut[26]), .S(n1078), .Q(n700) );
  MUX21X1 U1206 ( .IN1(\regfile[10][26] ), .IN2(AluOut[26]), .S(n1079), .Q(
        n699) );
  MUX21X1 U1207 ( .IN1(\regfile[11][26] ), .IN2(AluOut[26]), .S(n1080), .Q(
        n698) );
  MUX21X1 U1208 ( .IN1(\regfile[12][26] ), .IN2(AluOut[26]), .S(n1081), .Q(
        n697) );
  MUX21X1 U1209 ( .IN1(\regfile[13][26] ), .IN2(AluOut[26]), .S(n1082), .Q(
        n696) );
  MUX21X1 U1210 ( .IN1(\regfile[14][26] ), .IN2(AluOut[26]), .S(n1083), .Q(
        n695) );
  MUX21X1 U1211 ( .IN1(\regfile[15][26] ), .IN2(AluOut[26]), .S(n1084), .Q(
        n694) );
  AO221X1 U1212 ( .IN1(n1061), .IN2(AluOut[25]), .IN3(N181), .IN4(n1062), 
        .IN5(n1105), .Q(n693) );
  AO21X1 U1213 ( .IN1(IFID_A[25]), .IN2(n802), .IN3(n1106), .Q(n1105) );
  MUX21X1 U1214 ( .IN1(n1107), .IN2(n1108), .S(IFID_B[25]), .Q(n1106) );
  AO21X1 U1215 ( .IN1(IFID_A[25]), .IN2(n1067), .IN3(n802), .Q(n1108) );
  NOR2X0 U1216 ( .IN1(IFID_A[25]), .IN2(n1068), .QN(n1107) );
  MUX21X1 U1217 ( .IN1(\regfile[0][25] ), .IN2(AluOut[25]), .S(n1069), .Q(n692) );
  MUX21X1 U1218 ( .IN1(\regfile[1][25] ), .IN2(AluOut[25]), .S(n1070), .Q(n691) );
  MUX21X1 U1219 ( .IN1(\regfile[2][25] ), .IN2(AluOut[25]), .S(n1071), .Q(n690) );
  MUX21X1 U1220 ( .IN1(\regfile[3][25] ), .IN2(AluOut[25]), .S(n1072), .Q(n689) );
  MUX21X1 U1221 ( .IN1(\regfile[4][25] ), .IN2(AluOut[25]), .S(n1073), .Q(n688) );
  MUX21X1 U1222 ( .IN1(\regfile[5][25] ), .IN2(AluOut[25]), .S(n1074), .Q(n687) );
  MUX21X1 U1223 ( .IN1(\regfile[6][25] ), .IN2(AluOut[25]), .S(n1075), .Q(n686) );
  MUX21X1 U1224 ( .IN1(\regfile[7][25] ), .IN2(AluOut[25]), .S(n1076), .Q(n685) );
  MUX21X1 U1225 ( .IN1(\regfile[8][25] ), .IN2(AluOut[25]), .S(n1077), .Q(n684) );
  MUX21X1 U1226 ( .IN1(\regfile[9][25] ), .IN2(AluOut[25]), .S(n1078), .Q(n683) );
  MUX21X1 U1227 ( .IN1(\regfile[10][25] ), .IN2(AluOut[25]), .S(n1079), .Q(
        n682) );
  MUX21X1 U1228 ( .IN1(\regfile[11][25] ), .IN2(AluOut[25]), .S(n1080), .Q(
        n681) );
  MUX21X1 U1229 ( .IN1(\regfile[12][25] ), .IN2(AluOut[25]), .S(n1081), .Q(
        n680) );
  MUX21X1 U1230 ( .IN1(\regfile[13][25] ), .IN2(AluOut[25]), .S(n1082), .Q(
        n679) );
  MUX21X1 U1231 ( .IN1(\regfile[14][25] ), .IN2(AluOut[25]), .S(n1083), .Q(
        n678) );
  MUX21X1 U1232 ( .IN1(\regfile[15][25] ), .IN2(AluOut[25]), .S(n1084), .Q(
        n677) );
  AO221X1 U1233 ( .IN1(n1061), .IN2(AluOut[24]), .IN3(N180), .IN4(n1062), 
        .IN5(n1109), .Q(n676) );
  AO21X1 U1234 ( .IN1(IFID_A[24]), .IN2(n801), .IN3(n1110), .Q(n1109) );
  MUX21X1 U1235 ( .IN1(n1111), .IN2(n1112), .S(IFID_B[24]), .Q(n1110) );
  AO21X1 U1236 ( .IN1(IFID_A[24]), .IN2(n1067), .IN3(n801), .Q(n1112) );
  NOR2X0 U1237 ( .IN1(IFID_A[24]), .IN2(n1068), .QN(n1111) );
  MUX21X1 U1238 ( .IN1(\regfile[0][24] ), .IN2(AluOut[24]), .S(n1069), .Q(n675) );
  MUX21X1 U1239 ( .IN1(\regfile[1][24] ), .IN2(AluOut[24]), .S(n1070), .Q(n674) );
  MUX21X1 U1240 ( .IN1(\regfile[2][24] ), .IN2(AluOut[24]), .S(n1071), .Q(n673) );
  MUX21X1 U1241 ( .IN1(\regfile[3][24] ), .IN2(AluOut[24]), .S(n1072), .Q(n672) );
  MUX21X1 U1242 ( .IN1(\regfile[4][24] ), .IN2(AluOut[24]), .S(n1073), .Q(n671) );
  MUX21X1 U1243 ( .IN1(\regfile[5][24] ), .IN2(AluOut[24]), .S(n1074), .Q(n670) );
  MUX21X1 U1244 ( .IN1(\regfile[6][24] ), .IN2(AluOut[24]), .S(n1075), .Q(n669) );
  MUX21X1 U1245 ( .IN1(\regfile[7][24] ), .IN2(AluOut[24]), .S(n1076), .Q(n668) );
  MUX21X1 U1246 ( .IN1(\regfile[8][24] ), .IN2(AluOut[24]), .S(n1077), .Q(n667) );
  MUX21X1 U1247 ( .IN1(\regfile[9][24] ), .IN2(AluOut[24]), .S(n1078), .Q(n666) );
  MUX21X1 U1248 ( .IN1(\regfile[10][24] ), .IN2(AluOut[24]), .S(n1079), .Q(
        n665) );
  MUX21X1 U1249 ( .IN1(\regfile[11][24] ), .IN2(AluOut[24]), .S(n1080), .Q(
        n664) );
  MUX21X1 U1250 ( .IN1(\regfile[12][24] ), .IN2(AluOut[24]), .S(n1081), .Q(
        n663) );
  MUX21X1 U1251 ( .IN1(\regfile[13][24] ), .IN2(AluOut[24]), .S(n1082), .Q(
        n662) );
  MUX21X1 U1252 ( .IN1(\regfile[14][24] ), .IN2(AluOut[24]), .S(n1083), .Q(
        n661) );
  MUX21X1 U1253 ( .IN1(\regfile[15][24] ), .IN2(AluOut[24]), .S(n1084), .Q(
        n660) );
  AO221X1 U1254 ( .IN1(n1061), .IN2(AluOut[23]), .IN3(N179), .IN4(n1062), 
        .IN5(n1113), .Q(n659) );
  AO21X1 U1255 ( .IN1(IFID_A[23]), .IN2(n804), .IN3(n1114), .Q(n1113) );
  MUX21X1 U1256 ( .IN1(n1115), .IN2(n1116), .S(IFID_B[23]), .Q(n1114) );
  AO21X1 U1257 ( .IN1(IFID_A[23]), .IN2(n1067), .IN3(n804), .Q(n1116) );
  NOR2X0 U1258 ( .IN1(IFID_A[23]), .IN2(n1068), .QN(n1115) );
  MUX21X1 U1259 ( .IN1(\regfile[0][23] ), .IN2(AluOut[23]), .S(n1069), .Q(n658) );
  MUX21X1 U1260 ( .IN1(\regfile[1][23] ), .IN2(AluOut[23]), .S(n1070), .Q(n657) );
  MUX21X1 U1261 ( .IN1(\regfile[2][23] ), .IN2(AluOut[23]), .S(n1071), .Q(n656) );
  MUX21X1 U1262 ( .IN1(\regfile[3][23] ), .IN2(AluOut[23]), .S(n1072), .Q(n655) );
  MUX21X1 U1263 ( .IN1(\regfile[4][23] ), .IN2(AluOut[23]), .S(n1073), .Q(n654) );
  MUX21X1 U1264 ( .IN1(\regfile[5][23] ), .IN2(AluOut[23]), .S(n1074), .Q(n653) );
  MUX21X1 U1265 ( .IN1(\regfile[6][23] ), .IN2(AluOut[23]), .S(n1075), .Q(n652) );
  MUX21X1 U1266 ( .IN1(\regfile[7][23] ), .IN2(AluOut[23]), .S(n1076), .Q(n651) );
  MUX21X1 U1267 ( .IN1(\regfile[8][23] ), .IN2(AluOut[23]), .S(n1077), .Q(n650) );
  MUX21X1 U1268 ( .IN1(\regfile[9][23] ), .IN2(AluOut[23]), .S(n1078), .Q(n649) );
  MUX21X1 U1269 ( .IN1(\regfile[10][23] ), .IN2(AluOut[23]), .S(n1079), .Q(
        n648) );
  MUX21X1 U1270 ( .IN1(\regfile[11][23] ), .IN2(AluOut[23]), .S(n1080), .Q(
        n647) );
  MUX21X1 U1271 ( .IN1(\regfile[12][23] ), .IN2(AluOut[23]), .S(n1081), .Q(
        n646) );
  MUX21X1 U1272 ( .IN1(\regfile[13][23] ), .IN2(AluOut[23]), .S(n1082), .Q(
        n645) );
  MUX21X1 U1273 ( .IN1(\regfile[14][23] ), .IN2(AluOut[23]), .S(n1083), .Q(
        n644) );
  MUX21X1 U1274 ( .IN1(\regfile[15][23] ), .IN2(AluOut[23]), .S(n1084), .Q(
        n643) );
  AO221X1 U1275 ( .IN1(n1061), .IN2(AluOut[22]), .IN3(N178), .IN4(n1062), 
        .IN5(n1117), .Q(n642) );
  AO21X1 U1276 ( .IN1(IFID_A[22]), .IN2(n803), .IN3(n1118), .Q(n1117) );
  MUX21X1 U1277 ( .IN1(n1119), .IN2(n1120), .S(IFID_B[22]), .Q(n1118) );
  AO21X1 U1278 ( .IN1(IFID_A[22]), .IN2(n1067), .IN3(n803), .Q(n1120) );
  NOR2X0 U1279 ( .IN1(IFID_A[22]), .IN2(n1068), .QN(n1119) );
  MUX21X1 U1280 ( .IN1(\regfile[0][22] ), .IN2(AluOut[22]), .S(n1069), .Q(n641) );
  MUX21X1 U1281 ( .IN1(\regfile[1][22] ), .IN2(AluOut[22]), .S(n1070), .Q(n640) );
  MUX21X1 U1282 ( .IN1(\regfile[2][22] ), .IN2(AluOut[22]), .S(n1071), .Q(n639) );
  MUX21X1 U1283 ( .IN1(\regfile[3][22] ), .IN2(AluOut[22]), .S(n1072), .Q(n638) );
  MUX21X1 U1284 ( .IN1(\regfile[4][22] ), .IN2(AluOut[22]), .S(n1073), .Q(n637) );
  MUX21X1 U1285 ( .IN1(\regfile[5][22] ), .IN2(AluOut[22]), .S(n1074), .Q(n636) );
  MUX21X1 U1286 ( .IN1(\regfile[6][22] ), .IN2(AluOut[22]), .S(n1075), .Q(n635) );
  MUX21X1 U1287 ( .IN1(\regfile[7][22] ), .IN2(AluOut[22]), .S(n1076), .Q(n634) );
  MUX21X1 U1288 ( .IN1(\regfile[8][22] ), .IN2(AluOut[22]), .S(n1077), .Q(n633) );
  MUX21X1 U1289 ( .IN1(\regfile[9][22] ), .IN2(AluOut[22]), .S(n1078), .Q(n632) );
  MUX21X1 U1290 ( .IN1(\regfile[10][22] ), .IN2(AluOut[22]), .S(n1079), .Q(
        n631) );
  MUX21X1 U1291 ( .IN1(\regfile[11][22] ), .IN2(AluOut[22]), .S(n1080), .Q(
        n630) );
  MUX21X1 U1292 ( .IN1(\regfile[12][22] ), .IN2(AluOut[22]), .S(n1081), .Q(
        n629) );
  MUX21X1 U1293 ( .IN1(\regfile[13][22] ), .IN2(AluOut[22]), .S(n1082), .Q(
        n628) );
  MUX21X1 U1294 ( .IN1(\regfile[14][22] ), .IN2(AluOut[22]), .S(n1083), .Q(
        n627) );
  MUX21X1 U1295 ( .IN1(\regfile[15][22] ), .IN2(AluOut[22]), .S(n1084), .Q(
        n626) );
  AO221X1 U1296 ( .IN1(n1061), .IN2(AluOut[21]), .IN3(N177), .IN4(n1062), 
        .IN5(n1121), .Q(n625) );
  AO21X1 U1297 ( .IN1(IFID_A[21]), .IN2(n802), .IN3(n1122), .Q(n1121) );
  MUX21X1 U1298 ( .IN1(n1123), .IN2(n1124), .S(IFID_B[21]), .Q(n1122) );
  AO21X1 U1299 ( .IN1(IFID_A[21]), .IN2(n1067), .IN3(n802), .Q(n1124) );
  NOR2X0 U1300 ( .IN1(IFID_A[21]), .IN2(n1068), .QN(n1123) );
  MUX21X1 U1301 ( .IN1(\regfile[0][21] ), .IN2(AluOut[21]), .S(n1069), .Q(n624) );
  MUX21X1 U1302 ( .IN1(\regfile[1][21] ), .IN2(AluOut[21]), .S(n1070), .Q(n623) );
  MUX21X1 U1303 ( .IN1(\regfile[2][21] ), .IN2(AluOut[21]), .S(n1071), .Q(n622) );
  MUX21X1 U1304 ( .IN1(\regfile[3][21] ), .IN2(AluOut[21]), .S(n1072), .Q(n621) );
  MUX21X1 U1305 ( .IN1(\regfile[4][21] ), .IN2(AluOut[21]), .S(n1073), .Q(n620) );
  MUX21X1 U1306 ( .IN1(\regfile[5][21] ), .IN2(AluOut[21]), .S(n1074), .Q(n619) );
  MUX21X1 U1307 ( .IN1(\regfile[6][21] ), .IN2(AluOut[21]), .S(n1075), .Q(n618) );
  MUX21X1 U1308 ( .IN1(\regfile[7][21] ), .IN2(AluOut[21]), .S(n1076), .Q(n617) );
  MUX21X1 U1309 ( .IN1(\regfile[8][21] ), .IN2(AluOut[21]), .S(n1077), .Q(n616) );
  MUX21X1 U1310 ( .IN1(\regfile[9][21] ), .IN2(AluOut[21]), .S(n1078), .Q(n615) );
  MUX21X1 U1311 ( .IN1(\regfile[10][21] ), .IN2(AluOut[21]), .S(n1079), .Q(
        n614) );
  MUX21X1 U1312 ( .IN1(\regfile[11][21] ), .IN2(AluOut[21]), .S(n1080), .Q(
        n613) );
  MUX21X1 U1313 ( .IN1(\regfile[12][21] ), .IN2(AluOut[21]), .S(n1081), .Q(
        n612) );
  MUX21X1 U1314 ( .IN1(\regfile[13][21] ), .IN2(AluOut[21]), .S(n1082), .Q(
        n611) );
  MUX21X1 U1315 ( .IN1(\regfile[14][21] ), .IN2(AluOut[21]), .S(n1083), .Q(
        n610) );
  MUX21X1 U1316 ( .IN1(\regfile[15][21] ), .IN2(AluOut[21]), .S(n1084), .Q(
        n609) );
  AO221X1 U1317 ( .IN1(n1061), .IN2(AluOut[20]), .IN3(N176), .IN4(n1062), 
        .IN5(n1125), .Q(n608) );
  AO21X1 U1318 ( .IN1(IFID_A[20]), .IN2(n801), .IN3(n1126), .Q(n1125) );
  MUX21X1 U1319 ( .IN1(n1127), .IN2(n1128), .S(IFID_B[20]), .Q(n1126) );
  AO21X1 U1320 ( .IN1(IFID_A[20]), .IN2(n1067), .IN3(n801), .Q(n1128) );
  NOR2X0 U1321 ( .IN1(IFID_A[20]), .IN2(n1068), .QN(n1127) );
  MUX21X1 U1322 ( .IN1(\regfile[0][20] ), .IN2(AluOut[20]), .S(n1069), .Q(n607) );
  MUX21X1 U1323 ( .IN1(\regfile[1][20] ), .IN2(AluOut[20]), .S(n1070), .Q(n606) );
  MUX21X1 U1324 ( .IN1(\regfile[2][20] ), .IN2(AluOut[20]), .S(n1071), .Q(n605) );
  MUX21X1 U1325 ( .IN1(\regfile[3][20] ), .IN2(AluOut[20]), .S(n1072), .Q(n604) );
  MUX21X1 U1326 ( .IN1(\regfile[4][20] ), .IN2(AluOut[20]), .S(n1073), .Q(n603) );
  MUX21X1 U1327 ( .IN1(\regfile[5][20] ), .IN2(AluOut[20]), .S(n1074), .Q(n602) );
  MUX21X1 U1328 ( .IN1(\regfile[6][20] ), .IN2(AluOut[20]), .S(n1075), .Q(n601) );
  MUX21X1 U1329 ( .IN1(\regfile[7][20] ), .IN2(AluOut[20]), .S(n1076), .Q(n600) );
  MUX21X1 U1330 ( .IN1(\regfile[8][20] ), .IN2(AluOut[20]), .S(n1077), .Q(n599) );
  MUX21X1 U1331 ( .IN1(\regfile[9][20] ), .IN2(AluOut[20]), .S(n1078), .Q(n598) );
  MUX21X1 U1332 ( .IN1(\regfile[10][20] ), .IN2(AluOut[20]), .S(n1079), .Q(
        n597) );
  MUX21X1 U1333 ( .IN1(\regfile[11][20] ), .IN2(AluOut[20]), .S(n1080), .Q(
        n596) );
  MUX21X1 U1334 ( .IN1(\regfile[12][20] ), .IN2(AluOut[20]), .S(n1081), .Q(
        n595) );
  MUX21X1 U1335 ( .IN1(\regfile[13][20] ), .IN2(AluOut[20]), .S(n1082), .Q(
        n594) );
  MUX21X1 U1336 ( .IN1(\regfile[14][20] ), .IN2(AluOut[20]), .S(n1083), .Q(
        n593) );
  MUX21X1 U1337 ( .IN1(\regfile[15][20] ), .IN2(AluOut[20]), .S(n1084), .Q(
        n592) );
  AO221X1 U1338 ( .IN1(n1061), .IN2(AluOut[19]), .IN3(N175), .IN4(n1062), 
        .IN5(n1129), .Q(n591) );
  AO21X1 U1339 ( .IN1(IFID_A[19]), .IN2(n804), .IN3(n1130), .Q(n1129) );
  MUX21X1 U1340 ( .IN1(n1131), .IN2(n1132), .S(IFID_B[19]), .Q(n1130) );
  AO21X1 U1341 ( .IN1(IFID_A[19]), .IN2(n1067), .IN3(n804), .Q(n1132) );
  NOR2X0 U1342 ( .IN1(IFID_A[19]), .IN2(n1068), .QN(n1131) );
  MUX21X1 U1343 ( .IN1(\regfile[0][19] ), .IN2(AluOut[19]), .S(n1069), .Q(n590) );
  MUX21X1 U1344 ( .IN1(\regfile[1][19] ), .IN2(AluOut[19]), .S(n1070), .Q(n589) );
  MUX21X1 U1345 ( .IN1(\regfile[2][19] ), .IN2(AluOut[19]), .S(n1071), .Q(n588) );
  MUX21X1 U1346 ( .IN1(\regfile[3][19] ), .IN2(AluOut[19]), .S(n1072), .Q(n587) );
  MUX21X1 U1347 ( .IN1(\regfile[4][19] ), .IN2(AluOut[19]), .S(n1073), .Q(n586) );
  MUX21X1 U1348 ( .IN1(\regfile[5][19] ), .IN2(AluOut[19]), .S(n1074), .Q(n585) );
  MUX21X1 U1349 ( .IN1(\regfile[6][19] ), .IN2(AluOut[19]), .S(n1075), .Q(n584) );
  MUX21X1 U1350 ( .IN1(\regfile[7][19] ), .IN2(AluOut[19]), .S(n1076), .Q(n583) );
  MUX21X1 U1351 ( .IN1(\regfile[8][19] ), .IN2(AluOut[19]), .S(n1077), .Q(n582) );
  MUX21X1 U1352 ( .IN1(\regfile[9][19] ), .IN2(AluOut[19]), .S(n1078), .Q(n581) );
  MUX21X1 U1353 ( .IN1(\regfile[10][19] ), .IN2(AluOut[19]), .S(n1079), .Q(
        n580) );
  MUX21X1 U1354 ( .IN1(\regfile[11][19] ), .IN2(AluOut[19]), .S(n1080), .Q(
        n579) );
  MUX21X1 U1355 ( .IN1(\regfile[12][19] ), .IN2(AluOut[19]), .S(n1081), .Q(
        n578) );
  MUX21X1 U1356 ( .IN1(\regfile[13][19] ), .IN2(AluOut[19]), .S(n1082), .Q(
        n577) );
  MUX21X1 U1357 ( .IN1(\regfile[14][19] ), .IN2(AluOut[19]), .S(n1083), .Q(
        n576) );
  MUX21X1 U1358 ( .IN1(\regfile[15][19] ), .IN2(AluOut[19]), .S(n1084), .Q(
        n575) );
  AO221X1 U1359 ( .IN1(n1061), .IN2(AluOut[18]), .IN3(N174), .IN4(n1062), 
        .IN5(n1133), .Q(n574) );
  AO21X1 U1360 ( .IN1(IFID_A[18]), .IN2(n803), .IN3(n1134), .Q(n1133) );
  MUX21X1 U1361 ( .IN1(n1135), .IN2(n1136), .S(IFID_B[18]), .Q(n1134) );
  AO21X1 U1362 ( .IN1(IFID_A[18]), .IN2(n1067), .IN3(n803), .Q(n1136) );
  NOR2X0 U1363 ( .IN1(IFID_A[18]), .IN2(n1068), .QN(n1135) );
  MUX21X1 U1364 ( .IN1(\regfile[0][18] ), .IN2(AluOut[18]), .S(n1069), .Q(n573) );
  MUX21X1 U1365 ( .IN1(\regfile[1][18] ), .IN2(AluOut[18]), .S(n1070), .Q(n572) );
  MUX21X1 U1366 ( .IN1(\regfile[2][18] ), .IN2(AluOut[18]), .S(n1071), .Q(n571) );
  MUX21X1 U1367 ( .IN1(\regfile[3][18] ), .IN2(AluOut[18]), .S(n1072), .Q(n570) );
  MUX21X1 U1368 ( .IN1(\regfile[4][18] ), .IN2(AluOut[18]), .S(n1073), .Q(n569) );
  MUX21X1 U1369 ( .IN1(\regfile[5][18] ), .IN2(AluOut[18]), .S(n1074), .Q(n568) );
  MUX21X1 U1370 ( .IN1(\regfile[6][18] ), .IN2(AluOut[18]), .S(n1075), .Q(n567) );
  MUX21X1 U1371 ( .IN1(\regfile[7][18] ), .IN2(AluOut[18]), .S(n1076), .Q(n566) );
  MUX21X1 U1372 ( .IN1(\regfile[8][18] ), .IN2(AluOut[18]), .S(n1077), .Q(n565) );
  MUX21X1 U1373 ( .IN1(\regfile[9][18] ), .IN2(AluOut[18]), .S(n1078), .Q(n564) );
  MUX21X1 U1374 ( .IN1(\regfile[10][18] ), .IN2(AluOut[18]), .S(n1079), .Q(
        n563) );
  MUX21X1 U1375 ( .IN1(\regfile[11][18] ), .IN2(AluOut[18]), .S(n1080), .Q(
        n562) );
  MUX21X1 U1376 ( .IN1(\regfile[12][18] ), .IN2(AluOut[18]), .S(n1081), .Q(
        n561) );
  MUX21X1 U1377 ( .IN1(\regfile[13][18] ), .IN2(AluOut[18]), .S(n1082), .Q(
        n560) );
  MUX21X1 U1378 ( .IN1(\regfile[14][18] ), .IN2(AluOut[18]), .S(n1083), .Q(
        n559) );
  MUX21X1 U1379 ( .IN1(\regfile[15][18] ), .IN2(AluOut[18]), .S(n1084), .Q(
        n558) );
  AO221X1 U1380 ( .IN1(n1061), .IN2(AluOut[17]), .IN3(N173), .IN4(n1062), 
        .IN5(n1137), .Q(n557) );
  AO21X1 U1381 ( .IN1(IFID_A[17]), .IN2(n802), .IN3(n1138), .Q(n1137) );
  MUX21X1 U1382 ( .IN1(n1139), .IN2(n1140), .S(IFID_B[17]), .Q(n1138) );
  AO21X1 U1383 ( .IN1(IFID_A[17]), .IN2(n1067), .IN3(n802), .Q(n1140) );
  NOR2X0 U1384 ( .IN1(IFID_A[17]), .IN2(n1068), .QN(n1139) );
  MUX21X1 U1385 ( .IN1(\regfile[0][17] ), .IN2(AluOut[17]), .S(n1069), .Q(n556) );
  MUX21X1 U1386 ( .IN1(\regfile[1][17] ), .IN2(AluOut[17]), .S(n1070), .Q(n555) );
  MUX21X1 U1387 ( .IN1(\regfile[2][17] ), .IN2(AluOut[17]), .S(n1071), .Q(n554) );
  MUX21X1 U1388 ( .IN1(\regfile[3][17] ), .IN2(AluOut[17]), .S(n1072), .Q(n553) );
  MUX21X1 U1389 ( .IN1(\regfile[4][17] ), .IN2(AluOut[17]), .S(n1073), .Q(n552) );
  MUX21X1 U1390 ( .IN1(\regfile[5][17] ), .IN2(AluOut[17]), .S(n1074), .Q(n551) );
  MUX21X1 U1391 ( .IN1(\regfile[6][17] ), .IN2(AluOut[17]), .S(n1075), .Q(n550) );
  MUX21X1 U1392 ( .IN1(\regfile[7][17] ), .IN2(AluOut[17]), .S(n1076), .Q(n549) );
  MUX21X1 U1393 ( .IN1(\regfile[8][17] ), .IN2(AluOut[17]), .S(n1077), .Q(n548) );
  MUX21X1 U1394 ( .IN1(\regfile[9][17] ), .IN2(AluOut[17]), .S(n1078), .Q(n547) );
  MUX21X1 U1395 ( .IN1(\regfile[10][17] ), .IN2(AluOut[17]), .S(n1079), .Q(
        n546) );
  MUX21X1 U1396 ( .IN1(\regfile[11][17] ), .IN2(AluOut[17]), .S(n1080), .Q(
        n545) );
  MUX21X1 U1397 ( .IN1(\regfile[12][17] ), .IN2(AluOut[17]), .S(n1081), .Q(
        n544) );
  MUX21X1 U1398 ( .IN1(\regfile[13][17] ), .IN2(AluOut[17]), .S(n1082), .Q(
        n543) );
  MUX21X1 U1399 ( .IN1(\regfile[14][17] ), .IN2(AluOut[17]), .S(n1083), .Q(
        n542) );
  MUX21X1 U1400 ( .IN1(\regfile[15][17] ), .IN2(AluOut[17]), .S(n1084), .Q(
        n541) );
  AO221X1 U1401 ( .IN1(n1061), .IN2(AluOut[16]), .IN3(N172), .IN4(n1062), 
        .IN5(n1141), .Q(n540) );
  AO21X1 U1402 ( .IN1(IFID_A[16]), .IN2(n801), .IN3(n1142), .Q(n1141) );
  MUX21X1 U1403 ( .IN1(n1143), .IN2(n1144), .S(IFID_B[16]), .Q(n1142) );
  AO21X1 U1404 ( .IN1(IFID_A[16]), .IN2(n1067), .IN3(n801), .Q(n1144) );
  NOR2X0 U1405 ( .IN1(IFID_A[16]), .IN2(n1068), .QN(n1143) );
  MUX21X1 U1406 ( .IN1(\regfile[0][16] ), .IN2(AluOut[16]), .S(n1069), .Q(n539) );
  MUX21X1 U1407 ( .IN1(\regfile[1][16] ), .IN2(AluOut[16]), .S(n1070), .Q(n538) );
  MUX21X1 U1408 ( .IN1(\regfile[2][16] ), .IN2(AluOut[16]), .S(n1071), .Q(n537) );
  MUX21X1 U1409 ( .IN1(\regfile[3][16] ), .IN2(AluOut[16]), .S(n1072), .Q(n536) );
  MUX21X1 U1410 ( .IN1(\regfile[4][16] ), .IN2(AluOut[16]), .S(n1073), .Q(n535) );
  MUX21X1 U1411 ( .IN1(\regfile[5][16] ), .IN2(AluOut[16]), .S(n1074), .Q(n534) );
  MUX21X1 U1412 ( .IN1(\regfile[6][16] ), .IN2(AluOut[16]), .S(n1075), .Q(n533) );
  MUX21X1 U1413 ( .IN1(\regfile[7][16] ), .IN2(AluOut[16]), .S(n1076), .Q(n532) );
  MUX21X1 U1414 ( .IN1(\regfile[8][16] ), .IN2(AluOut[16]), .S(n1077), .Q(n531) );
  MUX21X1 U1415 ( .IN1(\regfile[9][16] ), .IN2(AluOut[16]), .S(n1078), .Q(n530) );
  MUX21X1 U1416 ( .IN1(\regfile[10][16] ), .IN2(AluOut[16]), .S(n1079), .Q(
        n529) );
  MUX21X1 U1417 ( .IN1(\regfile[11][16] ), .IN2(AluOut[16]), .S(n1080), .Q(
        n528) );
  MUX21X1 U1418 ( .IN1(\regfile[12][16] ), .IN2(AluOut[16]), .S(n1081), .Q(
        n527) );
  MUX21X1 U1419 ( .IN1(\regfile[13][16] ), .IN2(AluOut[16]), .S(n1082), .Q(
        n526) );
  MUX21X1 U1420 ( .IN1(\regfile[14][16] ), .IN2(AluOut[16]), .S(n1083), .Q(
        n525) );
  MUX21X1 U1421 ( .IN1(\regfile[15][16] ), .IN2(AluOut[16]), .S(n1084), .Q(
        n524) );
  AO221X1 U1422 ( .IN1(n1061), .IN2(AluOut[15]), .IN3(N171), .IN4(n1062), 
        .IN5(n1145), .Q(n523) );
  AO21X1 U1423 ( .IN1(IFID_A[15]), .IN2(n804), .IN3(n1146), .Q(n1145) );
  MUX21X1 U1424 ( .IN1(n1147), .IN2(n1148), .S(IFID_B[15]), .Q(n1146) );
  AO21X1 U1425 ( .IN1(IFID_A[15]), .IN2(n1067), .IN3(n804), .Q(n1148) );
  NOR2X0 U1426 ( .IN1(IFID_A[15]), .IN2(n1068), .QN(n1147) );
  MUX21X1 U1427 ( .IN1(\regfile[0][15] ), .IN2(AluOut[15]), .S(n1069), .Q(n522) );
  MUX21X1 U1428 ( .IN1(\regfile[1][15] ), .IN2(AluOut[15]), .S(n1070), .Q(n521) );
  MUX21X1 U1429 ( .IN1(\regfile[2][15] ), .IN2(AluOut[15]), .S(n1071), .Q(n520) );
  MUX21X1 U1430 ( .IN1(\regfile[3][15] ), .IN2(AluOut[15]), .S(n1072), .Q(n519) );
  MUX21X1 U1431 ( .IN1(\regfile[4][15] ), .IN2(AluOut[15]), .S(n1073), .Q(n518) );
  MUX21X1 U1432 ( .IN1(\regfile[5][15] ), .IN2(AluOut[15]), .S(n1074), .Q(n517) );
  MUX21X1 U1433 ( .IN1(\regfile[6][15] ), .IN2(AluOut[15]), .S(n1075), .Q(n516) );
  MUX21X1 U1434 ( .IN1(\regfile[7][15] ), .IN2(AluOut[15]), .S(n1076), .Q(n515) );
  MUX21X1 U1435 ( .IN1(\regfile[8][15] ), .IN2(AluOut[15]), .S(n1077), .Q(n514) );
  MUX21X1 U1436 ( .IN1(\regfile[9][15] ), .IN2(AluOut[15]), .S(n1078), .Q(n513) );
  MUX21X1 U1437 ( .IN1(\regfile[10][15] ), .IN2(AluOut[15]), .S(n1079), .Q(
        n512) );
  MUX21X1 U1438 ( .IN1(\regfile[11][15] ), .IN2(AluOut[15]), .S(n1080), .Q(
        n511) );
  MUX21X1 U1439 ( .IN1(\regfile[12][15] ), .IN2(AluOut[15]), .S(n1081), .Q(
        n510) );
  MUX21X1 U1440 ( .IN1(\regfile[13][15] ), .IN2(AluOut[15]), .S(n1082), .Q(
        n509) );
  MUX21X1 U1441 ( .IN1(\regfile[14][15] ), .IN2(AluOut[15]), .S(n1083), .Q(
        n508) );
  MUX21X1 U1442 ( .IN1(\regfile[15][15] ), .IN2(AluOut[15]), .S(n1084), .Q(
        n507) );
  AO221X1 U1443 ( .IN1(n1061), .IN2(AluOut[14]), .IN3(N170), .IN4(n1062), 
        .IN5(n1149), .Q(n506) );
  AO21X1 U1444 ( .IN1(IFID_A[14]), .IN2(n803), .IN3(n1150), .Q(n1149) );
  MUX21X1 U1445 ( .IN1(n1151), .IN2(n1152), .S(IFID_B[14]), .Q(n1150) );
  AO21X1 U1446 ( .IN1(IFID_A[14]), .IN2(n1067), .IN3(n803), .Q(n1152) );
  NOR2X0 U1447 ( .IN1(IFID_A[14]), .IN2(n1068), .QN(n1151) );
  MUX21X1 U1448 ( .IN1(\regfile[0][14] ), .IN2(AluOut[14]), .S(n1069), .Q(n505) );
  MUX21X1 U1449 ( .IN1(\regfile[1][14] ), .IN2(AluOut[14]), .S(n1070), .Q(n504) );
  MUX21X1 U1450 ( .IN1(\regfile[2][14] ), .IN2(AluOut[14]), .S(n1071), .Q(n503) );
  MUX21X1 U1451 ( .IN1(\regfile[3][14] ), .IN2(AluOut[14]), .S(n1072), .Q(n502) );
  MUX21X1 U1452 ( .IN1(\regfile[4][14] ), .IN2(AluOut[14]), .S(n1073), .Q(n501) );
  MUX21X1 U1453 ( .IN1(\regfile[5][14] ), .IN2(AluOut[14]), .S(n1074), .Q(n500) );
  MUX21X1 U1454 ( .IN1(\regfile[6][14] ), .IN2(AluOut[14]), .S(n1075), .Q(n499) );
  MUX21X1 U1455 ( .IN1(\regfile[7][14] ), .IN2(AluOut[14]), .S(n1076), .Q(n498) );
  MUX21X1 U1456 ( .IN1(\regfile[8][14] ), .IN2(AluOut[14]), .S(n1077), .Q(n497) );
  MUX21X1 U1457 ( .IN1(\regfile[9][14] ), .IN2(AluOut[14]), .S(n1078), .Q(n496) );
  MUX21X1 U1458 ( .IN1(\regfile[10][14] ), .IN2(AluOut[14]), .S(n1079), .Q(
        n495) );
  MUX21X1 U1459 ( .IN1(\regfile[11][14] ), .IN2(AluOut[14]), .S(n1080), .Q(
        n494) );
  MUX21X1 U1460 ( .IN1(\regfile[12][14] ), .IN2(AluOut[14]), .S(n1081), .Q(
        n493) );
  MUX21X1 U1461 ( .IN1(\regfile[13][14] ), .IN2(AluOut[14]), .S(n1082), .Q(
        n492) );
  MUX21X1 U1462 ( .IN1(\regfile[14][14] ), .IN2(AluOut[14]), .S(n1083), .Q(
        n491) );
  MUX21X1 U1463 ( .IN1(\regfile[15][14] ), .IN2(AluOut[14]), .S(n1084), .Q(
        n490) );
  AO221X1 U1464 ( .IN1(n1061), .IN2(AluOut[13]), .IN3(N169), .IN4(n1062), 
        .IN5(n1153), .Q(n489) );
  AO21X1 U1465 ( .IN1(IFID_A[13]), .IN2(n802), .IN3(n1154), .Q(n1153) );
  MUX21X1 U1466 ( .IN1(n1155), .IN2(n1156), .S(IFID_B[13]), .Q(n1154) );
  AO21X1 U1467 ( .IN1(IFID_A[13]), .IN2(n1067), .IN3(n802), .Q(n1156) );
  NOR2X0 U1468 ( .IN1(IFID_A[13]), .IN2(n1068), .QN(n1155) );
  MUX21X1 U1469 ( .IN1(\regfile[0][13] ), .IN2(AluOut[13]), .S(n1069), .Q(n488) );
  MUX21X1 U1470 ( .IN1(\regfile[1][13] ), .IN2(AluOut[13]), .S(n1070), .Q(n487) );
  MUX21X1 U1471 ( .IN1(\regfile[2][13] ), .IN2(AluOut[13]), .S(n1071), .Q(n486) );
  MUX21X1 U1472 ( .IN1(\regfile[3][13] ), .IN2(AluOut[13]), .S(n1072), .Q(n485) );
  MUX21X1 U1473 ( .IN1(\regfile[4][13] ), .IN2(AluOut[13]), .S(n1073), .Q(n484) );
  MUX21X1 U1474 ( .IN1(\regfile[5][13] ), .IN2(AluOut[13]), .S(n1074), .Q(n483) );
  MUX21X1 U1475 ( .IN1(\regfile[6][13] ), .IN2(AluOut[13]), .S(n1075), .Q(n482) );
  MUX21X1 U1476 ( .IN1(\regfile[7][13] ), .IN2(AluOut[13]), .S(n1076), .Q(n481) );
  MUX21X1 U1477 ( .IN1(\regfile[8][13] ), .IN2(AluOut[13]), .S(n1077), .Q(n480) );
  MUX21X1 U1478 ( .IN1(\regfile[9][13] ), .IN2(AluOut[13]), .S(n1078), .Q(n479) );
  MUX21X1 U1479 ( .IN1(\regfile[10][13] ), .IN2(AluOut[13]), .S(n1079), .Q(
        n478) );
  MUX21X1 U1480 ( .IN1(\regfile[11][13] ), .IN2(AluOut[13]), .S(n1080), .Q(
        n477) );
  MUX21X1 U1481 ( .IN1(\regfile[12][13] ), .IN2(AluOut[13]), .S(n1081), .Q(
        n476) );
  MUX21X1 U1482 ( .IN1(\regfile[13][13] ), .IN2(AluOut[13]), .S(n1082), .Q(
        n475) );
  MUX21X1 U1483 ( .IN1(\regfile[14][13] ), .IN2(AluOut[13]), .S(n1083), .Q(
        n474) );
  MUX21X1 U1484 ( .IN1(\regfile[15][13] ), .IN2(AluOut[13]), .S(n1084), .Q(
        n473) );
  AO221X1 U1485 ( .IN1(n1061), .IN2(AluOut[12]), .IN3(N168), .IN4(n1062), 
        .IN5(n1157), .Q(n472) );
  AO21X1 U1486 ( .IN1(IFID_A[12]), .IN2(n801), .IN3(n1158), .Q(n1157) );
  MUX21X1 U1487 ( .IN1(n1159), .IN2(n1160), .S(IFID_B[12]), .Q(n1158) );
  AO21X1 U1488 ( .IN1(IFID_A[12]), .IN2(n1067), .IN3(n801), .Q(n1160) );
  NOR2X0 U1489 ( .IN1(IFID_A[12]), .IN2(n1068), .QN(n1159) );
  MUX21X1 U1490 ( .IN1(\regfile[0][12] ), .IN2(AluOut[12]), .S(n1069), .Q(n471) );
  MUX21X1 U1491 ( .IN1(\regfile[1][12] ), .IN2(AluOut[12]), .S(n1070), .Q(n470) );
  MUX21X1 U1492 ( .IN1(\regfile[2][12] ), .IN2(AluOut[12]), .S(n1071), .Q(n469) );
  MUX21X1 U1493 ( .IN1(\regfile[3][12] ), .IN2(AluOut[12]), .S(n1072), .Q(n468) );
  MUX21X1 U1494 ( .IN1(\regfile[4][12] ), .IN2(AluOut[12]), .S(n1073), .Q(n467) );
  MUX21X1 U1495 ( .IN1(\regfile[5][12] ), .IN2(AluOut[12]), .S(n1074), .Q(n466) );
  MUX21X1 U1496 ( .IN1(\regfile[6][12] ), .IN2(AluOut[12]), .S(n1075), .Q(n465) );
  MUX21X1 U1497 ( .IN1(\regfile[7][12] ), .IN2(AluOut[12]), .S(n1076), .Q(n464) );
  MUX21X1 U1498 ( .IN1(\regfile[8][12] ), .IN2(AluOut[12]), .S(n1077), .Q(n463) );
  MUX21X1 U1499 ( .IN1(\regfile[9][12] ), .IN2(AluOut[12]), .S(n1078), .Q(n462) );
  MUX21X1 U1500 ( .IN1(\regfile[10][12] ), .IN2(AluOut[12]), .S(n1079), .Q(
        n461) );
  MUX21X1 U1501 ( .IN1(\regfile[11][12] ), .IN2(AluOut[12]), .S(n1080), .Q(
        n460) );
  MUX21X1 U1502 ( .IN1(\regfile[12][12] ), .IN2(AluOut[12]), .S(n1081), .Q(
        n459) );
  MUX21X1 U1503 ( .IN1(\regfile[13][12] ), .IN2(AluOut[12]), .S(n1082), .Q(
        n458) );
  MUX21X1 U1504 ( .IN1(\regfile[14][12] ), .IN2(AluOut[12]), .S(n1083), .Q(
        n457) );
  MUX21X1 U1505 ( .IN1(\regfile[15][12] ), .IN2(AluOut[12]), .S(n1084), .Q(
        n456) );
  AO221X1 U1506 ( .IN1(n1061), .IN2(AluOut[11]), .IN3(N167), .IN4(n1062), 
        .IN5(n1161), .Q(n455) );
  AO21X1 U1507 ( .IN1(IFID_A[11]), .IN2(n804), .IN3(n1162), .Q(n1161) );
  MUX21X1 U1508 ( .IN1(n1163), .IN2(n1164), .S(IFID_B[11]), .Q(n1162) );
  AO21X1 U1509 ( .IN1(IFID_A[11]), .IN2(n1067), .IN3(n804), .Q(n1164) );
  NOR2X0 U1510 ( .IN1(IFID_A[11]), .IN2(n1068), .QN(n1163) );
  MUX21X1 U1511 ( .IN1(\regfile[0][11] ), .IN2(AluOut[11]), .S(n1069), .Q(n454) );
  MUX21X1 U1512 ( .IN1(\regfile[1][11] ), .IN2(AluOut[11]), .S(n1070), .Q(n453) );
  MUX21X1 U1513 ( .IN1(\regfile[2][11] ), .IN2(AluOut[11]), .S(n1071), .Q(n452) );
  MUX21X1 U1514 ( .IN1(\regfile[3][11] ), .IN2(AluOut[11]), .S(n1072), .Q(n451) );
  MUX21X1 U1515 ( .IN1(\regfile[4][11] ), .IN2(AluOut[11]), .S(n1073), .Q(n450) );
  MUX21X1 U1516 ( .IN1(\regfile[5][11] ), .IN2(AluOut[11]), .S(n1074), .Q(n449) );
  MUX21X1 U1517 ( .IN1(\regfile[6][11] ), .IN2(AluOut[11]), .S(n1075), .Q(n448) );
  MUX21X1 U1518 ( .IN1(\regfile[7][11] ), .IN2(AluOut[11]), .S(n1076), .Q(n447) );
  MUX21X1 U1519 ( .IN1(\regfile[8][11] ), .IN2(AluOut[11]), .S(n1077), .Q(n446) );
  MUX21X1 U1520 ( .IN1(\regfile[9][11] ), .IN2(AluOut[11]), .S(n1078), .Q(n445) );
  MUX21X1 U1521 ( .IN1(\regfile[10][11] ), .IN2(AluOut[11]), .S(n1079), .Q(
        n444) );
  MUX21X1 U1522 ( .IN1(\regfile[11][11] ), .IN2(AluOut[11]), .S(n1080), .Q(
        n443) );
  MUX21X1 U1523 ( .IN1(\regfile[12][11] ), .IN2(AluOut[11]), .S(n1081), .Q(
        n442) );
  MUX21X1 U1524 ( .IN1(\regfile[13][11] ), .IN2(AluOut[11]), .S(n1082), .Q(
        n441) );
  MUX21X1 U1525 ( .IN1(\regfile[14][11] ), .IN2(AluOut[11]), .S(n1083), .Q(
        n440) );
  MUX21X1 U1526 ( .IN1(\regfile[15][11] ), .IN2(AluOut[11]), .S(n1084), .Q(
        n439) );
  AO221X1 U1527 ( .IN1(n1061), .IN2(AluOut[10]), .IN3(N166), .IN4(n1062), 
        .IN5(n1165), .Q(n438) );
  AO21X1 U1528 ( .IN1(IFID_A[10]), .IN2(n803), .IN3(n1166), .Q(n1165) );
  MUX21X1 U1529 ( .IN1(n1167), .IN2(n1168), .S(IFID_B[10]), .Q(n1166) );
  AO21X1 U1530 ( .IN1(IFID_A[10]), .IN2(n1067), .IN3(n803), .Q(n1168) );
  NOR2X0 U1531 ( .IN1(IFID_A[10]), .IN2(n1068), .QN(n1167) );
  MUX21X1 U1532 ( .IN1(\regfile[0][10] ), .IN2(AluOut[10]), .S(n1069), .Q(n437) );
  MUX21X1 U1533 ( .IN1(\regfile[1][10] ), .IN2(AluOut[10]), .S(n1070), .Q(n436) );
  MUX21X1 U1534 ( .IN1(\regfile[2][10] ), .IN2(AluOut[10]), .S(n1071), .Q(n435) );
  MUX21X1 U1535 ( .IN1(\regfile[3][10] ), .IN2(AluOut[10]), .S(n1072), .Q(n434) );
  MUX21X1 U1536 ( .IN1(\regfile[4][10] ), .IN2(AluOut[10]), .S(n1073), .Q(n433) );
  MUX21X1 U1537 ( .IN1(\regfile[5][10] ), .IN2(AluOut[10]), .S(n1074), .Q(n432) );
  MUX21X1 U1538 ( .IN1(\regfile[6][10] ), .IN2(AluOut[10]), .S(n1075), .Q(n431) );
  MUX21X1 U1539 ( .IN1(\regfile[7][10] ), .IN2(AluOut[10]), .S(n1076), .Q(n430) );
  MUX21X1 U1540 ( .IN1(\regfile[8][10] ), .IN2(AluOut[10]), .S(n1077), .Q(n429) );
  MUX21X1 U1541 ( .IN1(\regfile[9][10] ), .IN2(AluOut[10]), .S(n1078), .Q(n428) );
  MUX21X1 U1542 ( .IN1(\regfile[10][10] ), .IN2(AluOut[10]), .S(n1079), .Q(
        n427) );
  MUX21X1 U1543 ( .IN1(\regfile[11][10] ), .IN2(AluOut[10]), .S(n1080), .Q(
        n426) );
  MUX21X1 U1544 ( .IN1(\regfile[12][10] ), .IN2(AluOut[10]), .S(n1081), .Q(
        n425) );
  MUX21X1 U1545 ( .IN1(\regfile[13][10] ), .IN2(AluOut[10]), .S(n1082), .Q(
        n424) );
  MUX21X1 U1546 ( .IN1(\regfile[14][10] ), .IN2(AluOut[10]), .S(n1083), .Q(
        n423) );
  MUX21X1 U1547 ( .IN1(\regfile[15][10] ), .IN2(AluOut[10]), .S(n1084), .Q(
        n422) );
  AO221X1 U1548 ( .IN1(n1061), .IN2(AluOut[9]), .IN3(N165), .IN4(n1062), .IN5(
        n1169), .Q(n421) );
  AO21X1 U1549 ( .IN1(IFID_A[9]), .IN2(n802), .IN3(n1170), .Q(n1169) );
  MUX21X1 U1550 ( .IN1(n1171), .IN2(n1172), .S(IFID_B[9]), .Q(n1170) );
  AO21X1 U1551 ( .IN1(IFID_A[9]), .IN2(n1067), .IN3(n802), .Q(n1172) );
  NOR2X0 U1552 ( .IN1(IFID_A[9]), .IN2(n1068), .QN(n1171) );
  MUX21X1 U1553 ( .IN1(\regfile[0][9] ), .IN2(AluOut[9]), .S(n1069), .Q(n420)
         );
  MUX21X1 U1554 ( .IN1(\regfile[1][9] ), .IN2(AluOut[9]), .S(n1070), .Q(n419)
         );
  MUX21X1 U1555 ( .IN1(\regfile[2][9] ), .IN2(AluOut[9]), .S(n1071), .Q(n418)
         );
  MUX21X1 U1556 ( .IN1(\regfile[3][9] ), .IN2(AluOut[9]), .S(n1072), .Q(n417)
         );
  MUX21X1 U1557 ( .IN1(\regfile[4][9] ), .IN2(AluOut[9]), .S(n1073), .Q(n416)
         );
  MUX21X1 U1558 ( .IN1(\regfile[5][9] ), .IN2(AluOut[9]), .S(n1074), .Q(n415)
         );
  MUX21X1 U1559 ( .IN1(\regfile[6][9] ), .IN2(AluOut[9]), .S(n1075), .Q(n414)
         );
  MUX21X1 U1560 ( .IN1(\regfile[7][9] ), .IN2(AluOut[9]), .S(n1076), .Q(n413)
         );
  MUX21X1 U1561 ( .IN1(\regfile[8][9] ), .IN2(AluOut[9]), .S(n1077), .Q(n412)
         );
  MUX21X1 U1562 ( .IN1(\regfile[9][9] ), .IN2(AluOut[9]), .S(n1078), .Q(n411)
         );
  MUX21X1 U1563 ( .IN1(\regfile[10][9] ), .IN2(AluOut[9]), .S(n1079), .Q(n410)
         );
  MUX21X1 U1564 ( .IN1(\regfile[11][9] ), .IN2(AluOut[9]), .S(n1080), .Q(n409)
         );
  MUX21X1 U1565 ( .IN1(\regfile[12][9] ), .IN2(AluOut[9]), .S(n1081), .Q(n408)
         );
  MUX21X1 U1566 ( .IN1(\regfile[13][9] ), .IN2(AluOut[9]), .S(n1082), .Q(n407)
         );
  MUX21X1 U1567 ( .IN1(\regfile[14][9] ), .IN2(AluOut[9]), .S(n1083), .Q(n406)
         );
  MUX21X1 U1568 ( .IN1(\regfile[15][9] ), .IN2(AluOut[9]), .S(n1084), .Q(n405)
         );
  AO221X1 U1569 ( .IN1(n1061), .IN2(AluOut[8]), .IN3(N164), .IN4(n1062), .IN5(
        n1173), .Q(n404) );
  AO21X1 U1570 ( .IN1(IFID_A[8]), .IN2(n801), .IN3(n1174), .Q(n1173) );
  MUX21X1 U1571 ( .IN1(n1175), .IN2(n1176), .S(IFID_B[8]), .Q(n1174) );
  AO21X1 U1572 ( .IN1(IFID_A[8]), .IN2(n1067), .IN3(n801), .Q(n1176) );
  NOR2X0 U1573 ( .IN1(IFID_A[8]), .IN2(n1068), .QN(n1175) );
  MUX21X1 U1574 ( .IN1(\regfile[0][8] ), .IN2(AluOut[8]), .S(n1069), .Q(n403)
         );
  MUX21X1 U1575 ( .IN1(\regfile[1][8] ), .IN2(AluOut[8]), .S(n1070), .Q(n402)
         );
  MUX21X1 U1576 ( .IN1(\regfile[2][8] ), .IN2(AluOut[8]), .S(n1071), .Q(n401)
         );
  MUX21X1 U1577 ( .IN1(\regfile[3][8] ), .IN2(AluOut[8]), .S(n1072), .Q(n400)
         );
  MUX21X1 U1578 ( .IN1(\regfile[4][8] ), .IN2(AluOut[8]), .S(n1073), .Q(n399)
         );
  MUX21X1 U1579 ( .IN1(\regfile[5][8] ), .IN2(AluOut[8]), .S(n1074), .Q(n398)
         );
  MUX21X1 U1580 ( .IN1(\regfile[6][8] ), .IN2(AluOut[8]), .S(n1075), .Q(n397)
         );
  MUX21X1 U1581 ( .IN1(\regfile[7][8] ), .IN2(AluOut[8]), .S(n1076), .Q(n396)
         );
  MUX21X1 U1582 ( .IN1(\regfile[8][8] ), .IN2(AluOut[8]), .S(n1077), .Q(n395)
         );
  MUX21X1 U1583 ( .IN1(\regfile[9][8] ), .IN2(AluOut[8]), .S(n1078), .Q(n394)
         );
  MUX21X1 U1584 ( .IN1(\regfile[10][8] ), .IN2(AluOut[8]), .S(n1079), .Q(n393)
         );
  MUX21X1 U1585 ( .IN1(\regfile[11][8] ), .IN2(AluOut[8]), .S(n1080), .Q(n392)
         );
  MUX21X1 U1586 ( .IN1(\regfile[12][8] ), .IN2(AluOut[8]), .S(n1081), .Q(n391)
         );
  MUX21X1 U1587 ( .IN1(\regfile[13][8] ), .IN2(AluOut[8]), .S(n1082), .Q(n390)
         );
  MUX21X1 U1588 ( .IN1(\regfile[14][8] ), .IN2(AluOut[8]), .S(n1083), .Q(n389)
         );
  MUX21X1 U1589 ( .IN1(\regfile[15][8] ), .IN2(AluOut[8]), .S(n1084), .Q(n388)
         );
  AO221X1 U1590 ( .IN1(n1061), .IN2(AluOut[7]), .IN3(N163), .IN4(n1062), .IN5(
        n1177), .Q(n387) );
  AO21X1 U1591 ( .IN1(IFID_A[7]), .IN2(n804), .IN3(n1178), .Q(n1177) );
  MUX21X1 U1592 ( .IN1(n1179), .IN2(n1180), .S(IFID_B[7]), .Q(n1178) );
  AO21X1 U1593 ( .IN1(IFID_A[7]), .IN2(n1067), .IN3(n804), .Q(n1180) );
  NOR2X0 U1594 ( .IN1(IFID_A[7]), .IN2(n1068), .QN(n1179) );
  MUX21X1 U1595 ( .IN1(\regfile[0][7] ), .IN2(AluOut[7]), .S(n1069), .Q(n386)
         );
  MUX21X1 U1596 ( .IN1(\regfile[1][7] ), .IN2(AluOut[7]), .S(n1070), .Q(n385)
         );
  MUX21X1 U1597 ( .IN1(\regfile[2][7] ), .IN2(AluOut[7]), .S(n1071), .Q(n384)
         );
  MUX21X1 U1598 ( .IN1(\regfile[3][7] ), .IN2(AluOut[7]), .S(n1072), .Q(n383)
         );
  MUX21X1 U1599 ( .IN1(\regfile[4][7] ), .IN2(AluOut[7]), .S(n1073), .Q(n382)
         );
  MUX21X1 U1600 ( .IN1(\regfile[5][7] ), .IN2(AluOut[7]), .S(n1074), .Q(n381)
         );
  MUX21X1 U1601 ( .IN1(\regfile[6][7] ), .IN2(AluOut[7]), .S(n1075), .Q(n380)
         );
  MUX21X1 U1602 ( .IN1(\regfile[7][7] ), .IN2(AluOut[7]), .S(n1076), .Q(n379)
         );
  MUX21X1 U1603 ( .IN1(\regfile[8][7] ), .IN2(AluOut[7]), .S(n1077), .Q(n378)
         );
  MUX21X1 U1604 ( .IN1(\regfile[9][7] ), .IN2(AluOut[7]), .S(n1078), .Q(n377)
         );
  MUX21X1 U1605 ( .IN1(\regfile[10][7] ), .IN2(AluOut[7]), .S(n1079), .Q(n376)
         );
  MUX21X1 U1606 ( .IN1(\regfile[11][7] ), .IN2(AluOut[7]), .S(n1080), .Q(n375)
         );
  MUX21X1 U1607 ( .IN1(\regfile[12][7] ), .IN2(AluOut[7]), .S(n1081), .Q(n374)
         );
  MUX21X1 U1608 ( .IN1(\regfile[13][7] ), .IN2(AluOut[7]), .S(n1082), .Q(n373)
         );
  MUX21X1 U1609 ( .IN1(\regfile[14][7] ), .IN2(AluOut[7]), .S(n1083), .Q(n372)
         );
  MUX21X1 U1610 ( .IN1(\regfile[15][7] ), .IN2(AluOut[7]), .S(n1084), .Q(n371)
         );
  AO221X1 U1611 ( .IN1(n1061), .IN2(AluOut[6]), .IN3(N162), .IN4(n1062), .IN5(
        n1181), .Q(n370) );
  AO21X1 U1612 ( .IN1(IFID_A[6]), .IN2(n803), .IN3(n1182), .Q(n1181) );
  MUX21X1 U1613 ( .IN1(n1183), .IN2(n1184), .S(IFID_B[6]), .Q(n1182) );
  AO21X1 U1614 ( .IN1(IFID_A[6]), .IN2(n1067), .IN3(n803), .Q(n1184) );
  NOR2X0 U1615 ( .IN1(IFID_A[6]), .IN2(n1068), .QN(n1183) );
  MUX21X1 U1616 ( .IN1(\regfile[0][6] ), .IN2(AluOut[6]), .S(n1069), .Q(n369)
         );
  MUX21X1 U1617 ( .IN1(\regfile[1][6] ), .IN2(AluOut[6]), .S(n1070), .Q(n368)
         );
  MUX21X1 U1618 ( .IN1(\regfile[2][6] ), .IN2(AluOut[6]), .S(n1071), .Q(n367)
         );
  MUX21X1 U1619 ( .IN1(\regfile[3][6] ), .IN2(AluOut[6]), .S(n1072), .Q(n366)
         );
  MUX21X1 U1620 ( .IN1(\regfile[4][6] ), .IN2(AluOut[6]), .S(n1073), .Q(n365)
         );
  MUX21X1 U1621 ( .IN1(\regfile[5][6] ), .IN2(AluOut[6]), .S(n1074), .Q(n364)
         );
  MUX21X1 U1622 ( .IN1(\regfile[6][6] ), .IN2(AluOut[6]), .S(n1075), .Q(n363)
         );
  MUX21X1 U1623 ( .IN1(\regfile[7][6] ), .IN2(AluOut[6]), .S(n1076), .Q(n362)
         );
  MUX21X1 U1624 ( .IN1(\regfile[8][6] ), .IN2(AluOut[6]), .S(n1077), .Q(n361)
         );
  MUX21X1 U1625 ( .IN1(\regfile[9][6] ), .IN2(AluOut[6]), .S(n1078), .Q(n360)
         );
  MUX21X1 U1626 ( .IN1(\regfile[10][6] ), .IN2(AluOut[6]), .S(n1079), .Q(n359)
         );
  MUX21X1 U1627 ( .IN1(\regfile[11][6] ), .IN2(AluOut[6]), .S(n1080), .Q(n358)
         );
  MUX21X1 U1628 ( .IN1(\regfile[12][6] ), .IN2(AluOut[6]), .S(n1081), .Q(n357)
         );
  MUX21X1 U1629 ( .IN1(\regfile[13][6] ), .IN2(AluOut[6]), .S(n1082), .Q(n356)
         );
  MUX21X1 U1630 ( .IN1(\regfile[14][6] ), .IN2(AluOut[6]), .S(n1083), .Q(n355)
         );
  MUX21X1 U1631 ( .IN1(\regfile[15][6] ), .IN2(AluOut[6]), .S(n1084), .Q(n354)
         );
  AO221X1 U1632 ( .IN1(n1061), .IN2(AluOut[5]), .IN3(N161), .IN4(n1062), .IN5(
        n1185), .Q(n353) );
  AO21X1 U1633 ( .IN1(IFID_A[5]), .IN2(n802), .IN3(n1186), .Q(n1185) );
  MUX21X1 U1634 ( .IN1(n1187), .IN2(n1188), .S(IFID_B[5]), .Q(n1186) );
  AO21X1 U1635 ( .IN1(IFID_A[5]), .IN2(n1067), .IN3(n802), .Q(n1188) );
  NOR2X0 U1636 ( .IN1(IFID_A[5]), .IN2(n1068), .QN(n1187) );
  MUX21X1 U1637 ( .IN1(\regfile[0][5] ), .IN2(AluOut[5]), .S(n1069), .Q(n352)
         );
  MUX21X1 U1638 ( .IN1(\regfile[1][5] ), .IN2(AluOut[5]), .S(n1070), .Q(n351)
         );
  MUX21X1 U1639 ( .IN1(\regfile[2][5] ), .IN2(AluOut[5]), .S(n1071), .Q(n350)
         );
  MUX21X1 U1640 ( .IN1(\regfile[3][5] ), .IN2(AluOut[5]), .S(n1072), .Q(n349)
         );
  MUX21X1 U1641 ( .IN1(\regfile[4][5] ), .IN2(AluOut[5]), .S(n1073), .Q(n348)
         );
  MUX21X1 U1642 ( .IN1(\regfile[5][5] ), .IN2(AluOut[5]), .S(n1074), .Q(n347)
         );
  MUX21X1 U1643 ( .IN1(\regfile[6][5] ), .IN2(AluOut[5]), .S(n1075), .Q(n346)
         );
  MUX21X1 U1644 ( .IN1(\regfile[7][5] ), .IN2(AluOut[5]), .S(n1076), .Q(n345)
         );
  MUX21X1 U1645 ( .IN1(\regfile[8][5] ), .IN2(AluOut[5]), .S(n1077), .Q(n344)
         );
  MUX21X1 U1646 ( .IN1(\regfile[9][5] ), .IN2(AluOut[5]), .S(n1078), .Q(n343)
         );
  MUX21X1 U1647 ( .IN1(\regfile[10][5] ), .IN2(AluOut[5]), .S(n1079), .Q(n342)
         );
  MUX21X1 U1648 ( .IN1(\regfile[11][5] ), .IN2(AluOut[5]), .S(n1080), .Q(n341)
         );
  MUX21X1 U1649 ( .IN1(\regfile[12][5] ), .IN2(AluOut[5]), .S(n1081), .Q(n340)
         );
  MUX21X1 U1650 ( .IN1(\regfile[13][5] ), .IN2(AluOut[5]), .S(n1082), .Q(n339)
         );
  MUX21X1 U1651 ( .IN1(\regfile[14][5] ), .IN2(AluOut[5]), .S(n1083), .Q(n338)
         );
  MUX21X1 U1652 ( .IN1(\regfile[15][5] ), .IN2(AluOut[5]), .S(n1084), .Q(n337)
         );
  AO221X1 U1653 ( .IN1(n1061), .IN2(AluOut[4]), .IN3(N160), .IN4(n1062), .IN5(
        n1189), .Q(n336) );
  AO21X1 U1654 ( .IN1(IFID_A[4]), .IN2(n801), .IN3(n1190), .Q(n1189) );
  MUX21X1 U1655 ( .IN1(n1191), .IN2(n1192), .S(IFID_B[4]), .Q(n1190) );
  AO21X1 U1656 ( .IN1(IFID_A[4]), .IN2(n1067), .IN3(n801), .Q(n1192) );
  NOR2X0 U1657 ( .IN1(IFID_A[4]), .IN2(n1068), .QN(n1191) );
  MUX21X1 U1658 ( .IN1(\regfile[0][4] ), .IN2(AluOut[4]), .S(n1069), .Q(n335)
         );
  MUX21X1 U1659 ( .IN1(\regfile[1][4] ), .IN2(AluOut[4]), .S(n1070), .Q(n334)
         );
  MUX21X1 U1660 ( .IN1(\regfile[2][4] ), .IN2(AluOut[4]), .S(n1071), .Q(n333)
         );
  MUX21X1 U1661 ( .IN1(\regfile[3][4] ), .IN2(AluOut[4]), .S(n1072), .Q(n332)
         );
  MUX21X1 U1662 ( .IN1(\regfile[4][4] ), .IN2(AluOut[4]), .S(n1073), .Q(n331)
         );
  MUX21X1 U1663 ( .IN1(\regfile[5][4] ), .IN2(AluOut[4]), .S(n1074), .Q(n330)
         );
  MUX21X1 U1664 ( .IN1(\regfile[6][4] ), .IN2(AluOut[4]), .S(n1075), .Q(n329)
         );
  MUX21X1 U1665 ( .IN1(\regfile[7][4] ), .IN2(AluOut[4]), .S(n1076), .Q(n328)
         );
  MUX21X1 U1666 ( .IN1(\regfile[8][4] ), .IN2(AluOut[4]), .S(n1077), .Q(n327)
         );
  MUX21X1 U1667 ( .IN1(\regfile[9][4] ), .IN2(AluOut[4]), .S(n1078), .Q(n326)
         );
  MUX21X1 U1668 ( .IN1(\regfile[10][4] ), .IN2(AluOut[4]), .S(n1079), .Q(n325)
         );
  MUX21X1 U1669 ( .IN1(\regfile[11][4] ), .IN2(AluOut[4]), .S(n1080), .Q(n324)
         );
  MUX21X1 U1670 ( .IN1(\regfile[12][4] ), .IN2(AluOut[4]), .S(n1081), .Q(n323)
         );
  MUX21X1 U1671 ( .IN1(\regfile[13][4] ), .IN2(AluOut[4]), .S(n1082), .Q(n322)
         );
  MUX21X1 U1672 ( .IN1(\regfile[14][4] ), .IN2(AluOut[4]), .S(n1083), .Q(n321)
         );
  MUX21X1 U1673 ( .IN1(\regfile[15][4] ), .IN2(AluOut[4]), .S(n1084), .Q(n320)
         );
  AO221X1 U1674 ( .IN1(n1061), .IN2(AluOut[3]), .IN3(N159), .IN4(n1062), .IN5(
        n1193), .Q(n319) );
  AO21X1 U1675 ( .IN1(IFID_A[3]), .IN2(n804), .IN3(n1194), .Q(n1193) );
  MUX21X1 U1676 ( .IN1(n1195), .IN2(n1196), .S(IFID_B[3]), .Q(n1194) );
  AO21X1 U1677 ( .IN1(IFID_A[3]), .IN2(n1067), .IN3(n804), .Q(n1196) );
  NOR2X0 U1678 ( .IN1(IFID_A[3]), .IN2(n1068), .QN(n1195) );
  MUX21X1 U1679 ( .IN1(\regfile[0][3] ), .IN2(AluOut[3]), .S(n1069), .Q(n318)
         );
  MUX21X1 U1680 ( .IN1(\regfile[1][3] ), .IN2(AluOut[3]), .S(n1070), .Q(n317)
         );
  MUX21X1 U1681 ( .IN1(\regfile[2][3] ), .IN2(AluOut[3]), .S(n1071), .Q(n316)
         );
  MUX21X1 U1682 ( .IN1(\regfile[3][3] ), .IN2(AluOut[3]), .S(n1072), .Q(n315)
         );
  MUX21X1 U1683 ( .IN1(\regfile[4][3] ), .IN2(AluOut[3]), .S(n1073), .Q(n314)
         );
  MUX21X1 U1684 ( .IN1(\regfile[5][3] ), .IN2(AluOut[3]), .S(n1074), .Q(n313)
         );
  MUX21X1 U1685 ( .IN1(\regfile[6][3] ), .IN2(AluOut[3]), .S(n1075), .Q(n312)
         );
  MUX21X1 U1686 ( .IN1(\regfile[7][3] ), .IN2(AluOut[3]), .S(n1076), .Q(n311)
         );
  MUX21X1 U1687 ( .IN1(\regfile[8][3] ), .IN2(AluOut[3]), .S(n1077), .Q(n310)
         );
  MUX21X1 U1688 ( .IN1(\regfile[9][3] ), .IN2(AluOut[3]), .S(n1078), .Q(n309)
         );
  MUX21X1 U1689 ( .IN1(\regfile[10][3] ), .IN2(AluOut[3]), .S(n1079), .Q(n308)
         );
  MUX21X1 U1690 ( .IN1(\regfile[11][3] ), .IN2(AluOut[3]), .S(n1080), .Q(n307)
         );
  MUX21X1 U1691 ( .IN1(\regfile[12][3] ), .IN2(AluOut[3]), .S(n1081), .Q(n306)
         );
  MUX21X1 U1692 ( .IN1(\regfile[13][3] ), .IN2(AluOut[3]), .S(n1082), .Q(n305)
         );
  MUX21X1 U1693 ( .IN1(\regfile[14][3] ), .IN2(AluOut[3]), .S(n1083), .Q(n304)
         );
  MUX21X1 U1694 ( .IN1(\regfile[15][3] ), .IN2(AluOut[3]), .S(n1084), .Q(n303)
         );
  AO221X1 U1695 ( .IN1(n1061), .IN2(AluOut[2]), .IN3(N158), .IN4(n1062), .IN5(
        n1197), .Q(n302) );
  AO21X1 U1696 ( .IN1(IFID_A[2]), .IN2(n803), .IN3(n1198), .Q(n1197) );
  MUX21X1 U1697 ( .IN1(n1199), .IN2(n1200), .S(IFID_B[2]), .Q(n1198) );
  AO21X1 U1698 ( .IN1(IFID_A[2]), .IN2(n1067), .IN3(n803), .Q(n1200) );
  NOR2X0 U1699 ( .IN1(IFID_A[2]), .IN2(n1068), .QN(n1199) );
  MUX21X1 U1700 ( .IN1(\regfile[0][2] ), .IN2(AluOut[2]), .S(n1069), .Q(n301)
         );
  MUX21X1 U1701 ( .IN1(\regfile[1][2] ), .IN2(AluOut[2]), .S(n1070), .Q(n300)
         );
  MUX21X1 U1702 ( .IN1(\regfile[2][2] ), .IN2(AluOut[2]), .S(n1071), .Q(n299)
         );
  MUX21X1 U1703 ( .IN1(\regfile[3][2] ), .IN2(AluOut[2]), .S(n1072), .Q(n298)
         );
  MUX21X1 U1704 ( .IN1(\regfile[4][2] ), .IN2(AluOut[2]), .S(n1073), .Q(n297)
         );
  MUX21X1 U1705 ( .IN1(\regfile[5][2] ), .IN2(AluOut[2]), .S(n1074), .Q(n296)
         );
  MUX21X1 U1706 ( .IN1(\regfile[6][2] ), .IN2(AluOut[2]), .S(n1075), .Q(n295)
         );
  MUX21X1 U1707 ( .IN1(\regfile[7][2] ), .IN2(AluOut[2]), .S(n1076), .Q(n294)
         );
  MUX21X1 U1708 ( .IN1(\regfile[8][2] ), .IN2(AluOut[2]), .S(n1077), .Q(n293)
         );
  MUX21X1 U1709 ( .IN1(\regfile[9][2] ), .IN2(AluOut[2]), .S(n1078), .Q(n292)
         );
  MUX21X1 U1710 ( .IN1(\regfile[10][2] ), .IN2(AluOut[2]), .S(n1079), .Q(n291)
         );
  MUX21X1 U1711 ( .IN1(\regfile[11][2] ), .IN2(AluOut[2]), .S(n1080), .Q(n290)
         );
  MUX21X1 U1712 ( .IN1(\regfile[12][2] ), .IN2(AluOut[2]), .S(n1081), .Q(n289)
         );
  MUX21X1 U1713 ( .IN1(\regfile[13][2] ), .IN2(AluOut[2]), .S(n1082), .Q(n288)
         );
  MUX21X1 U1714 ( .IN1(\regfile[14][2] ), .IN2(AluOut[2]), .S(n1083), .Q(n287)
         );
  MUX21X1 U1715 ( .IN1(\regfile[15][2] ), .IN2(AluOut[2]), .S(n1084), .Q(n286)
         );
  AO221X1 U1716 ( .IN1(n1061), .IN2(AluOut[1]), .IN3(N157), .IN4(n1062), .IN5(
        n1201), .Q(n285) );
  AO21X1 U1717 ( .IN1(IFID_A[1]), .IN2(n802), .IN3(n1202), .Q(n1201) );
  MUX21X1 U1718 ( .IN1(n1203), .IN2(n1204), .S(IFID_B[1]), .Q(n1202) );
  AO21X1 U1719 ( .IN1(IFID_A[1]), .IN2(n1067), .IN3(n802), .Q(n1204) );
  NOR2X0 U1720 ( .IN1(IFID_A[1]), .IN2(n1068), .QN(n1203) );
  INVX0 U1721 ( .INP(n1205), .ZN(n1061) );
  MUX21X1 U1722 ( .IN1(\regfile[0][1] ), .IN2(AluOut[1]), .S(n1069), .Q(n284)
         );
  MUX21X1 U1723 ( .IN1(\regfile[1][1] ), .IN2(AluOut[1]), .S(n1070), .Q(n283)
         );
  MUX21X1 U1724 ( .IN1(\regfile[2][1] ), .IN2(AluOut[1]), .S(n1071), .Q(n282)
         );
  MUX21X1 U1725 ( .IN1(\regfile[3][1] ), .IN2(AluOut[1]), .S(n1072), .Q(n281)
         );
  MUX21X1 U1726 ( .IN1(\regfile[4][1] ), .IN2(AluOut[1]), .S(n1073), .Q(n280)
         );
  MUX21X1 U1727 ( .IN1(\regfile[5][1] ), .IN2(AluOut[1]), .S(n1074), .Q(n279)
         );
  MUX21X1 U1728 ( .IN1(\regfile[6][1] ), .IN2(AluOut[1]), .S(n1075), .Q(n278)
         );
  MUX21X1 U1729 ( .IN1(\regfile[7][1] ), .IN2(AluOut[1]), .S(n1076), .Q(n277)
         );
  MUX21X1 U1730 ( .IN1(\regfile[8][1] ), .IN2(AluOut[1]), .S(n1077), .Q(n276)
         );
  MUX21X1 U1731 ( .IN1(\regfile[9][1] ), .IN2(AluOut[1]), .S(n1078), .Q(n275)
         );
  MUX21X1 U1732 ( .IN1(\regfile[10][1] ), .IN2(AluOut[1]), .S(n1079), .Q(n274)
         );
  MUX21X1 U1733 ( .IN1(\regfile[11][1] ), .IN2(AluOut[1]), .S(n1080), .Q(n273)
         );
  MUX21X1 U1734 ( .IN1(\regfile[12][1] ), .IN2(AluOut[1]), .S(n1081), .Q(n272)
         );
  MUX21X1 U1735 ( .IN1(\regfile[13][1] ), .IN2(AluOut[1]), .S(n1082), .Q(n271)
         );
  MUX21X1 U1736 ( .IN1(\regfile[14][1] ), .IN2(AluOut[1]), .S(n1083), .Q(n270)
         );
  MUX21X1 U1737 ( .IN1(\regfile[15][1] ), .IN2(AluOut[1]), .S(n1084), .Q(n269)
         );
  NAND4X0 U1738 ( .IN1(n1206), .IN2(n1207), .IN3(n1208), .IN4(n1209), .QN(n268) );
  OA221X1 U1739 ( .IN1(n216), .IN2(n1205), .IN3(IFID_A[31]), .IN4(n1210), 
        .IN5(n1211), .Q(n1209) );
  AO22X1 U1740 ( .IN1(n1212), .IN2(n1213), .IN3(n1210), .IN4(n1214), .Q(n1211)
         );
  NAND3X0 U1741 ( .IN1(instr[12]), .IN2(n1215), .IN3(n1216), .QN(n1214) );
  AO221X1 U1742 ( .IN1(IFID_A[30]), .IN2(n1217), .IN3(IFID_A[29]), .IN4(n1218), 
        .IN5(n1219), .Q(n1213) );
  OA221X1 U1743 ( .IN1(IFID_A[29]), .IN2(n1218), .IN3(IFID_A[28]), .IN4(n1220), 
        .IN5(n1221), .Q(n1219) );
  AO221X1 U1744 ( .IN1(IFID_A[28]), .IN2(n1220), .IN3(IFID_A[27]), .IN4(n1222), 
        .IN5(n1223), .Q(n1221) );
  OA221X1 U1745 ( .IN1(IFID_A[27]), .IN2(n1222), .IN3(IFID_A[26]), .IN4(n1224), 
        .IN5(n1225), .Q(n1223) );
  AO221X1 U1746 ( .IN1(IFID_A[26]), .IN2(n1224), .IN3(IFID_A[25]), .IN4(n1226), 
        .IN5(n1227), .Q(n1225) );
  OA221X1 U1747 ( .IN1(IFID_A[25]), .IN2(n1226), .IN3(IFID_A[24]), .IN4(n1228), 
        .IN5(n1229), .Q(n1227) );
  AO221X1 U1748 ( .IN1(IFID_A[24]), .IN2(n1228), .IN3(IFID_A[23]), .IN4(n1230), 
        .IN5(n1231), .Q(n1229) );
  OA221X1 U1749 ( .IN1(IFID_A[23]), .IN2(n1230), .IN3(IFID_A[22]), .IN4(n1232), 
        .IN5(n1233), .Q(n1231) );
  AO221X1 U1750 ( .IN1(IFID_A[22]), .IN2(n1232), .IN3(IFID_A[21]), .IN4(n1234), 
        .IN5(n1235), .Q(n1233) );
  OA221X1 U1751 ( .IN1(IFID_A[21]), .IN2(n1234), .IN3(IFID_A[20]), .IN4(n1236), 
        .IN5(n1237), .Q(n1235) );
  AO221X1 U1752 ( .IN1(IFID_A[20]), .IN2(n1236), .IN3(IFID_A[19]), .IN4(n1238), 
        .IN5(n1239), .Q(n1237) );
  OA221X1 U1753 ( .IN1(IFID_A[19]), .IN2(n1238), .IN3(IFID_A[18]), .IN4(n1240), 
        .IN5(n1241), .Q(n1239) );
  AO221X1 U1754 ( .IN1(IFID_A[18]), .IN2(n1240), .IN3(IFID_A[17]), .IN4(n1242), 
        .IN5(n1243), .Q(n1241) );
  OA221X1 U1755 ( .IN1(IFID_A[17]), .IN2(n1242), .IN3(IFID_A[16]), .IN4(n1244), 
        .IN5(n1245), .Q(n1243) );
  AO221X1 U1756 ( .IN1(IFID_A[16]), .IN2(n1244), .IN3(IFID_A[15]), .IN4(n1246), 
        .IN5(n1247), .Q(n1245) );
  OA221X1 U1757 ( .IN1(IFID_A[15]), .IN2(n1246), .IN3(IFID_A[14]), .IN4(n1248), 
        .IN5(n1249), .Q(n1247) );
  AO221X1 U1758 ( .IN1(IFID_A[14]), .IN2(n1248), .IN3(IFID_A[13]), .IN4(n1250), 
        .IN5(n1251), .Q(n1249) );
  OA221X1 U1759 ( .IN1(IFID_A[13]), .IN2(n1250), .IN3(IFID_A[12]), .IN4(n1252), 
        .IN5(n1253), .Q(n1251) );
  AO221X1 U1760 ( .IN1(IFID_A[12]), .IN2(n1252), .IN3(IFID_A[11]), .IN4(n1254), 
        .IN5(n1255), .Q(n1253) );
  OA221X1 U1761 ( .IN1(IFID_A[11]), .IN2(n1254), .IN3(IFID_A[10]), .IN4(n1256), 
        .IN5(n1257), .Q(n1255) );
  AO221X1 U1762 ( .IN1(IFID_A[10]), .IN2(n1256), .IN3(IFID_A[9]), .IN4(n1258), 
        .IN5(n1259), .Q(n1257) );
  OA221X1 U1763 ( .IN1(IFID_A[9]), .IN2(n1258), .IN3(IFID_A[8]), .IN4(n1260), 
        .IN5(n1261), .Q(n1259) );
  AO221X1 U1764 ( .IN1(IFID_A[8]), .IN2(n1260), .IN3(IFID_A[7]), .IN4(n1262), 
        .IN5(n1263), .Q(n1261) );
  OA221X1 U1765 ( .IN1(IFID_A[7]), .IN2(n1262), .IN3(IFID_A[6]), .IN4(n1264), 
        .IN5(n1265), .Q(n1263) );
  AO221X1 U1766 ( .IN1(IFID_A[6]), .IN2(n1264), .IN3(IFID_A[5]), .IN4(n1266), 
        .IN5(n1267), .Q(n1265) );
  OA221X1 U1767 ( .IN1(IFID_A[5]), .IN2(n1266), .IN3(IFID_A[4]), .IN4(n1268), 
        .IN5(n1269), .Q(n1267) );
  AO221X1 U1768 ( .IN1(IFID_A[4]), .IN2(n1268), .IN3(IFID_A[3]), .IN4(n1270), 
        .IN5(n1271), .Q(n1269) );
  OA222X1 U1769 ( .IN1(IFID_A[3]), .IN2(n1270), .IN3(n1272), .IN4(n1273), 
        .IN5(IFID_A[2]), .IN6(n1274), .Q(n1271) );
  INVX0 U1770 ( .INP(IFID_B[2]), .ZN(n1273) );
  AND2X1 U1771 ( .IN1(IFID_A[2]), .IN2(n1274), .Q(n1272) );
  AOI22X1 U1772 ( .IN1(n1275), .IN2(n1276), .IN3(IFID_B[1]), .IN4(n1277), .QN(
        n1274) );
  OR2X1 U1773 ( .IN1(n1276), .IN2(n1275), .Q(n1277) );
  INVX0 U1774 ( .INP(IFID_A[1]), .ZN(n1276) );
  NOR2X0 U1775 ( .IN1(n1278), .IN2(IFID_A[0]), .QN(n1275) );
  INVX0 U1776 ( .INP(IFID_B[3]), .ZN(n1270) );
  INVX0 U1777 ( .INP(IFID_B[4]), .ZN(n1268) );
  INVX0 U1778 ( .INP(IFID_B[5]), .ZN(n1266) );
  INVX0 U1779 ( .INP(IFID_B[6]), .ZN(n1264) );
  INVX0 U1780 ( .INP(IFID_B[7]), .ZN(n1262) );
  INVX0 U1781 ( .INP(IFID_B[8]), .ZN(n1260) );
  INVX0 U1782 ( .INP(IFID_B[9]), .ZN(n1258) );
  INVX0 U1783 ( .INP(IFID_B[10]), .ZN(n1256) );
  INVX0 U1784 ( .INP(IFID_B[11]), .ZN(n1254) );
  INVX0 U1785 ( .INP(IFID_B[12]), .ZN(n1252) );
  INVX0 U1786 ( .INP(IFID_B[13]), .ZN(n1250) );
  INVX0 U1787 ( .INP(IFID_B[14]), .ZN(n1248) );
  INVX0 U1788 ( .INP(IFID_B[15]), .ZN(n1246) );
  INVX0 U1789 ( .INP(IFID_B[16]), .ZN(n1244) );
  INVX0 U1790 ( .INP(IFID_B[17]), .ZN(n1242) );
  INVX0 U1791 ( .INP(IFID_B[18]), .ZN(n1240) );
  INVX0 U1792 ( .INP(IFID_B[19]), .ZN(n1238) );
  INVX0 U1793 ( .INP(IFID_B[20]), .ZN(n1236) );
  INVX0 U1794 ( .INP(IFID_B[21]), .ZN(n1234) );
  INVX0 U1795 ( .INP(IFID_B[22]), .ZN(n1232) );
  INVX0 U1796 ( .INP(IFID_B[23]), .ZN(n1230) );
  INVX0 U1797 ( .INP(IFID_B[24]), .ZN(n1228) );
  INVX0 U1798 ( .INP(IFID_B[25]), .ZN(n1226) );
  INVX0 U1799 ( .INP(IFID_B[26]), .ZN(n1224) );
  INVX0 U1800 ( .INP(IFID_B[27]), .ZN(n1222) );
  INVX0 U1801 ( .INP(IFID_B[28]), .ZN(n1220) );
  INVX0 U1802 ( .INP(IFID_B[29]), .ZN(n1218) );
  OR2X1 U1803 ( .IN1(n1217), .IN2(IFID_A[30]), .Q(n1212) );
  INVX0 U1804 ( .INP(IFID_B[30]), .ZN(n1217) );
  NAND3X0 U1805 ( .IN1(IFID_B[31]), .IN2(instr[12]), .IN3(n1216), .QN(n1210)
         );
  INVX0 U1806 ( .INP(n1279), .ZN(n1216) );
  NAND4X0 U1807 ( .IN1(n1280), .IN2(n1068), .IN3(n1281), .IN4(n1279), .QN(
        n1205) );
  NAND3X0 U1808 ( .IN1(instr[13]), .IN2(n1282), .IN3(instr[14]), .QN(n1279) );
  MUX21X1 U1809 ( .IN1(n1283), .IN2(n1284), .S(n1278), .Q(n1208) );
  INVX0 U1810 ( .INP(IFID_B[0]), .ZN(n1278) );
  OR2X1 U1811 ( .IN1(n1068), .IN2(IFID_A[0]), .Q(n1284) );
  NAND4X0 U1812 ( .IN1(instr[15]), .IN2(instr[14]), .IN3(n1285), .IN4(n1286), 
        .QN(n1068) );
  AOI21X1 U1813 ( .IN1(n1067), .IN2(IFID_A[0]), .IN3(n801), .QN(n1283) );
  INVX0 U1814 ( .INP(n1280), .ZN(n1067) );
  NAND2X0 U1815 ( .IN1(N156), .IN2(n1062), .QN(n1207) );
  NAND2X0 U1816 ( .IN1(IFID_A[0]), .IN2(n804), .QN(n1206) );
  NAND3X0 U1817 ( .IN1(n1287), .IN2(n1282), .IN3(n1286), .QN(n1280) );
  INVX0 U1818 ( .INP(instr[13]), .ZN(n1286) );
  MUX21X1 U1819 ( .IN1(\regfile[0][0] ), .IN2(AluOut[0]), .S(n1069), .Q(n267)
         );
  AND2X1 U1820 ( .IN1(n1288), .IN2(n1289), .Q(n1069) );
  MUX21X1 U1821 ( .IN1(\regfile[1][0] ), .IN2(AluOut[0]), .S(n1070), .Q(n266)
         );
  AND2X1 U1822 ( .IN1(n1290), .IN2(n1289), .Q(n1070) );
  MUX21X1 U1823 ( .IN1(\regfile[2][0] ), .IN2(AluOut[0]), .S(n1071), .Q(n265)
         );
  AND2X1 U1824 ( .IN1(n1291), .IN2(n1288), .Q(n1071) );
  MUX21X1 U1825 ( .IN1(\regfile[3][0] ), .IN2(AluOut[0]), .S(n1072), .Q(n264)
         );
  AND2X1 U1826 ( .IN1(n1291), .IN2(n1290), .Q(n1072) );
  MUX21X1 U1827 ( .IN1(\regfile[4][0] ), .IN2(AluOut[0]), .S(n1073), .Q(n263)
         );
  AND2X1 U1828 ( .IN1(n1292), .IN2(n1289), .Q(n1073) );
  MUX21X1 U1829 ( .IN1(\regfile[5][0] ), .IN2(AluOut[0]), .S(n1074), .Q(n262)
         );
  AND2X1 U1830 ( .IN1(n1293), .IN2(n1289), .Q(n1074) );
  NOR2X0 U1831 ( .IN1(n1315), .IN2(n1316), .QN(n1289) );
  MUX21X1 U1832 ( .IN1(\regfile[6][0] ), .IN2(AluOut[0]), .S(n1075), .Q(n261)
         );
  AND2X1 U1833 ( .IN1(n1292), .IN2(n1291), .Q(n1075) );
  MUX21X1 U1834 ( .IN1(\regfile[7][0] ), .IN2(AluOut[0]), .S(n1076), .Q(n260)
         );
  AND2X1 U1835 ( .IN1(n1293), .IN2(n1291), .Q(n1076) );
  NOR2X0 U1836 ( .IN1(n799), .IN2(n1315), .QN(n1291) );
  MUX21X1 U1837 ( .IN1(\regfile[8][0] ), .IN2(AluOut[0]), .S(n1077), .Q(n259)
         );
  AND2X1 U1838 ( .IN1(n1294), .IN2(n1288), .Q(n1077) );
  MUX21X1 U1839 ( .IN1(\regfile[9][0] ), .IN2(AluOut[0]), .S(n1078), .Q(n258)
         );
  AND2X1 U1840 ( .IN1(n1294), .IN2(n1290), .Q(n1078) );
  MUX21X1 U1841 ( .IN1(\regfile[10][0] ), .IN2(AluOut[0]), .S(n1079), .Q(n257)
         );
  AND2X1 U1842 ( .IN1(n1295), .IN2(n1288), .Q(n1079) );
  NOR2X0 U1843 ( .IN1(n1313), .IN2(n1314), .QN(n1288) );
  MUX21X1 U1844 ( .IN1(\regfile[11][0] ), .IN2(AluOut[0]), .S(n1080), .Q(n256)
         );
  AND2X1 U1845 ( .IN1(n1295), .IN2(n1290), .Q(n1080) );
  NOR2X0 U1846 ( .IN1(n800), .IN2(n1313), .QN(n1290) );
  MUX21X1 U1847 ( .IN1(\regfile[12][0] ), .IN2(AluOut[0]), .S(n1081), .Q(n255)
         );
  AND2X1 U1848 ( .IN1(n1294), .IN2(n1292), .Q(n1081) );
  MUX21X1 U1849 ( .IN1(\regfile[13][0] ), .IN2(AluOut[0]), .S(n1082), .Q(n254)
         );
  AND2X1 U1850 ( .IN1(n1294), .IN2(n1293), .Q(n1082) );
  AND2X1 U1851 ( .IN1(n1315), .IN2(n799), .Q(n1294) );
  MUX21X1 U1852 ( .IN1(\regfile[14][0] ), .IN2(AluOut[0]), .S(n1083), .Q(n253)
         );
  AND2X1 U1853 ( .IN1(n1295), .IN2(n1292), .Q(n1083) );
  AND2X1 U1854 ( .IN1(n1313), .IN2(n800), .Q(n1292) );
  MUX21X1 U1855 ( .IN1(\regfile[15][0] ), .IN2(AluOut[0]), .S(n1084), .Q(n252)
         );
  AND2X1 U1856 ( .IN1(n1295), .IN2(n1293), .Q(n1084) );
  AND2X1 U1857 ( .IN1(n1313), .IN2(n1314), .Q(n1293) );
  AND2X1 U1858 ( .IN1(n1315), .IN2(n1316), .Q(n1295) );
  AND2X1 U1859 ( .IN1(n1296), .IN2(n1297), .Q(Zero) );
  NOR4X0 U1860 ( .IN1(n1298), .IN2(n1299), .IN3(n1300), .IN4(n1301), .QN(n1297) );
  NAND4X0 U1861 ( .IN1(n231), .IN2(n230), .IN3(n229), .IN4(n228), .QN(n1301)
         );
  NAND4X0 U1862 ( .IN1(n227), .IN2(n226), .IN3(n225), .IN4(n224), .QN(n1300)
         );
  NAND4X0 U1863 ( .IN1(n223), .IN2(n222), .IN3(n221), .IN4(n220), .QN(n1299)
         );
  NAND4X0 U1864 ( .IN1(n219), .IN2(n218), .IN3(n217), .IN4(n216), .QN(n1298)
         );
  NOR4X0 U1865 ( .IN1(n1302), .IN2(n1303), .IN3(n1304), .IN4(n1305), .QN(n1296) );
  NAND4X0 U1866 ( .IN1(n251), .IN2(n246), .IN3(n245), .IN4(n244), .QN(n1305)
         );
  NAND4X0 U1867 ( .IN1(n243), .IN2(n242), .IN3(n241), .IN4(n240), .QN(n1304)
         );
  NAND4X0 U1868 ( .IN1(n239), .IN2(n238), .IN3(n237), .IN4(n236), .QN(n1303)
         );
  NAND4X0 U1869 ( .IN1(n235), .IN2(n234), .IN3(n233), .IN4(n232), .QN(n1302)
         );
  MUX21X1 U1870 ( .IN1(n1306), .IN2(n1307), .S(N187), .Q(N257) );
  OAI21X1 U1871 ( .IN1(n1308), .IN2(n1309), .IN3(n1310), .QN(n1307) );
  NAND3X0 U1872 ( .IN1(n1311), .IN2(n1287), .IN3(n1062), .QN(n1310) );
  AOI21X1 U1873 ( .IN1(n1215), .IN2(IFID_B[31]), .IN3(N188), .QN(n1308) );
  AO22X1 U1874 ( .IN1(n1317), .IN2(n1287), .IN3(n1312), .IN4(n1318), .Q(n1306)
         );
  NAND2X0 U1875 ( .IN1(instr[14]), .IN2(n1062), .QN(n1309) );
  INVX0 U1876 ( .INP(n1281), .ZN(n1062) );
  NOR2X0 U1877 ( .IN1(IFID_B[31]), .IN2(n1215), .QN(n1312) );
  INVX0 U1878 ( .INP(IFID_A[31]), .ZN(n1215) );
  INVX0 U1879 ( .INP(instr[14]), .ZN(n1287) );
  NOR2X0 U1880 ( .IN1(n1311), .IN2(n1281), .QN(n1317) );
  NAND3X0 U1881 ( .IN1(n1285), .IN2(n1282), .IN3(instr[13]), .QN(n1281) );
  INVX0 U1882 ( .INP(instr[15]), .ZN(n1282) );
  INVX0 U1883 ( .INP(instr[12]), .ZN(n1285) );
  INVX0 U1884 ( .INP(N188), .ZN(n1311) );
endmodule



module thumb_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [33:0] carry;
  wire   [32:0] B_AS;
  assign B_AS[32] = ADD_SUB;

  FADDX1 U1_31 ( .A(A[31]), .B(B_AS[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B_AS[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B_AS[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B_AS[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B_AS[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B_AS[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B_AS[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B_AS[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B_AS[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B_AS[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B_AS[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B_AS[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B_AS[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B_AS[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B_AS[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B_AS[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B_AS[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FADDX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FADDX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FADDX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FADDX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FADDX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FADDX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FADDX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FADDX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0]) );
  XOR2X1 U1 ( .IN1(B_AS[32]), .IN2(carry[32]), .Q(SUM[32]) );
  XOR2X1 U2 ( .IN1(CI), .IN2(B_AS[32]), .Q(carry[0]) );
  XOR2X1 U3 ( .IN1(B[9]), .IN2(B_AS[32]), .Q(B_AS[9]) );
  XOR2X1 U4 ( .IN1(B[8]), .IN2(B_AS[32]), .Q(B_AS[8]) );
  XOR2X1 U5 ( .IN1(B[7]), .IN2(B_AS[32]), .Q(B_AS[7]) );
  XOR2X1 U6 ( .IN1(B[6]), .IN2(B_AS[32]), .Q(B_AS[6]) );
  XOR2X1 U7 ( .IN1(B[5]), .IN2(B_AS[32]), .Q(B_AS[5]) );
  XOR2X1 U8 ( .IN1(B[4]), .IN2(B_AS[32]), .Q(B_AS[4]) );
  XOR2X1 U9 ( .IN1(B[3]), .IN2(B_AS[32]), .Q(B_AS[3]) );
  XOR2X1 U10 ( .IN1(B[31]), .IN2(B_AS[32]), .Q(B_AS[31]) );
  XOR2X1 U11 ( .IN1(B[30]), .IN2(B_AS[32]), .Q(B_AS[30]) );
  XOR2X1 U12 ( .IN1(B[2]), .IN2(B_AS[32]), .Q(B_AS[2]) );
  XOR2X1 U13 ( .IN1(B[29]), .IN2(B_AS[32]), .Q(B_AS[29]) );
  XOR2X1 U14 ( .IN1(B[28]), .IN2(B_AS[32]), .Q(B_AS[28]) );
  XOR2X1 U15 ( .IN1(B[27]), .IN2(B_AS[32]), .Q(B_AS[27]) );
  XOR2X1 U16 ( .IN1(B[26]), .IN2(B_AS[32]), .Q(B_AS[26]) );
  XOR2X1 U17 ( .IN1(B[25]), .IN2(B_AS[32]), .Q(B_AS[25]) );
  XOR2X1 U18 ( .IN1(B[24]), .IN2(B_AS[32]), .Q(B_AS[24]) );
  XOR2X1 U19 ( .IN1(B[23]), .IN2(B_AS[32]), .Q(B_AS[23]) );
  XOR2X1 U20 ( .IN1(B[22]), .IN2(B_AS[32]), .Q(B_AS[22]) );
  XOR2X1 U21 ( .IN1(B[21]), .IN2(B_AS[32]), .Q(B_AS[21]) );
  XOR2X1 U22 ( .IN1(B[20]), .IN2(B_AS[32]), .Q(B_AS[20]) );
  XOR2X1 U23 ( .IN1(B[1]), .IN2(B_AS[32]), .Q(B_AS[1]) );
  XOR2X1 U24 ( .IN1(B[19]), .IN2(B_AS[32]), .Q(B_AS[19]) );
  XOR2X1 U25 ( .IN1(B[18]), .IN2(B_AS[32]), .Q(B_AS[18]) );
  XOR2X1 U26 ( .IN1(B[17]), .IN2(B_AS[32]), .Q(B_AS[17]) );
  XOR2X1 U27 ( .IN1(B[16]), .IN2(B_AS[32]), .Q(B_AS[16]) );
  XOR2X1 U28 ( .IN1(B[15]), .IN2(B_AS[32]), .Q(B_AS[15]) );
  XOR2X1 U29 ( .IN1(B[14]), .IN2(B_AS[32]), .Q(B_AS[14]) );
  XOR2X1 U30 ( .IN1(B[13]), .IN2(B_AS[32]), .Q(B_AS[13]) );
  XOR2X1 U31 ( .IN1(B[12]), .IN2(B_AS[32]), .Q(B_AS[12]) );
  XOR2X1 U32 ( .IN1(B[11]), .IN2(B_AS[32]), .Q(B_AS[11]) );
  XOR2X1 U33 ( .IN1(B[10]), .IN2(B_AS[32]), .Q(B_AS[10]) );
  XOR2X1 U34 ( .IN1(B[0]), .IN2(B_AS[32]), .Q(B_AS[0]) );
endmodule


module thumb_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [32:1] carry;
  assign SUM[1] = A[1];
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  AND2X1 U1 ( .IN1(A[2]), .IN2(B[2]), .Q(n1) );
  AND2X1 U2 ( .IN1(A[7]), .IN2(carry[7]), .Q(n2) );
  AND2X1 U3 ( .IN1(A[8]), .IN2(n2), .Q(n3) );
  AND2X1 U4 ( .IN1(A[9]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(A[10]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(A[11]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(A[12]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(A[13]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(A[14]), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(A[15]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(A[16]), .IN2(n10), .Q(n11) );
  AND2X1 U12 ( .IN1(A[17]), .IN2(n11), .Q(n12) );
  AND2X1 U13 ( .IN1(A[18]), .IN2(n12), .Q(n13) );
  AND2X1 U14 ( .IN1(A[19]), .IN2(n13), .Q(n14) );
  AND2X1 U15 ( .IN1(A[20]), .IN2(n14), .Q(n15) );
  AND2X1 U16 ( .IN1(A[21]), .IN2(n15), .Q(n16) );
  AND2X1 U17 ( .IN1(A[22]), .IN2(n16), .Q(n17) );
  AND2X1 U18 ( .IN1(A[23]), .IN2(n17), .Q(n18) );
  AND2X1 U19 ( .IN1(A[28]), .IN2(n25), .Q(n19) );
  AND2X1 U20 ( .IN1(A[24]), .IN2(n18), .Q(n20) );
  AND2X1 U21 ( .IN1(A[29]), .IN2(n19), .Q(n21) );
  AND2X1 U22 ( .IN1(A[25]), .IN2(n20), .Q(n22) );
  AND2X1 U23 ( .IN1(A[30]), .IN2(n21), .Q(n23) );
  AND2X1 U24 ( .IN1(A[26]), .IN2(n22), .Q(n24) );
  AND2X1 U25 ( .IN1(A[27]), .IN2(n24), .Q(n25) );
  AND2X1 U26 ( .IN1(A[31]), .IN2(n23), .Q(SUM[32]) );
  XOR2X1 U27 ( .IN1(A[31]), .IN2(n23), .Q(SUM[31]) );
  XOR2X1 U28 ( .IN1(A[30]), .IN2(n21), .Q(SUM[30]) );
  XOR2X1 U29 ( .IN1(A[29]), .IN2(n19), .Q(SUM[29]) );
  XOR2X1 U30 ( .IN1(A[28]), .IN2(n25), .Q(SUM[28]) );
  XOR2X1 U31 ( .IN1(A[27]), .IN2(n24), .Q(SUM[27]) );
  XOR2X1 U32 ( .IN1(A[26]), .IN2(n22), .Q(SUM[26]) );
  XOR2X1 U33 ( .IN1(A[25]), .IN2(n20), .Q(SUM[25]) );
  XOR2X1 U34 ( .IN1(A[24]), .IN2(n18), .Q(SUM[24]) );
  XOR2X1 U35 ( .IN1(A[23]), .IN2(n17), .Q(SUM[23]) );
  XOR2X1 U36 ( .IN1(A[22]), .IN2(n16), .Q(SUM[22]) );
  XOR2X1 U37 ( .IN1(A[21]), .IN2(n15), .Q(SUM[21]) );
  XOR2X1 U38 ( .IN1(A[20]), .IN2(n14), .Q(SUM[20]) );
  XOR2X1 U39 ( .IN1(A[19]), .IN2(n13), .Q(SUM[19]) );
  XOR2X1 U40 ( .IN1(A[18]), .IN2(n12), .Q(SUM[18]) );
  XOR2X1 U41 ( .IN1(A[17]), .IN2(n11), .Q(SUM[17]) );
  XOR2X1 U42 ( .IN1(A[16]), .IN2(n10), .Q(SUM[16]) );
  XOR2X1 U43 ( .IN1(A[15]), .IN2(n9), .Q(SUM[15]) );
  XOR2X1 U44 ( .IN1(A[14]), .IN2(n8), .Q(SUM[14]) );
  XOR2X1 U45 ( .IN1(A[13]), .IN2(n7), .Q(SUM[13]) );
  XOR2X1 U46 ( .IN1(A[12]), .IN2(n6), .Q(SUM[12]) );
  XOR2X1 U47 ( .IN1(A[11]), .IN2(n5), .Q(SUM[11]) );
  XOR2X1 U48 ( .IN1(A[10]), .IN2(n4), .Q(SUM[10]) );
  XOR2X1 U49 ( .IN1(A[9]), .IN2(n3), .Q(SUM[9]) );
  XOR2X1 U50 ( .IN1(A[8]), .IN2(n2), .Q(SUM[8]) );
  XOR2X1 U51 ( .IN1(A[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U52 ( .IN1(A[2]), .IN2(B[2]), .Q(SUM[2]) );
endmodule


module thumb_DW01_add_1 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23;
  wire   [32:1] carry;
  assign SUM[1] = A[1];
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(n2), .CO(carry[4]), .S(SUM[3]) );
  AND2X1 U1 ( .IN1(A[31]), .IN2(n23), .Q(SUM[32]) );
  AND2X1 U2 ( .IN1(A[2]), .IN2(B[2]), .Q(n2) );
  AND2X1 U3 ( .IN1(A[10]), .IN2(carry[10]), .Q(n3) );
  AND2X1 U4 ( .IN1(A[11]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(A[12]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(A[13]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(A[14]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(A[15]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(A[16]), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(A[17]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(A[18]), .IN2(n10), .Q(n11) );
  AND2X1 U12 ( .IN1(A[19]), .IN2(n11), .Q(n12) );
  AND2X1 U13 ( .IN1(A[20]), .IN2(n12), .Q(n13) );
  AND2X1 U14 ( .IN1(A[21]), .IN2(n13), .Q(n14) );
  AND2X1 U15 ( .IN1(A[22]), .IN2(n14), .Q(n15) );
  AND2X1 U16 ( .IN1(A[23]), .IN2(n15), .Q(n16) );
  AND2X1 U17 ( .IN1(A[24]), .IN2(n16), .Q(n17) );
  AND2X1 U18 ( .IN1(A[25]), .IN2(n17), .Q(n18) );
  AND2X1 U19 ( .IN1(A[26]), .IN2(n18), .Q(n19) );
  AND2X1 U20 ( .IN1(A[27]), .IN2(n19), .Q(n20) );
  AND2X1 U21 ( .IN1(A[28]), .IN2(n20), .Q(n21) );
  AND2X1 U22 ( .IN1(A[29]), .IN2(n21), .Q(n22) );
  AND2X1 U23 ( .IN1(A[30]), .IN2(n22), .Q(n23) );
  XOR2X1 U24 ( .IN1(A[31]), .IN2(n23), .Q(SUM[31]) );
  XOR2X1 U25 ( .IN1(A[30]), .IN2(n22), .Q(SUM[30]) );
  XOR2X1 U26 ( .IN1(A[29]), .IN2(n21), .Q(SUM[29]) );
  XOR2X1 U27 ( .IN1(A[28]), .IN2(n20), .Q(SUM[28]) );
  XOR2X1 U28 ( .IN1(A[27]), .IN2(n19), .Q(SUM[27]) );
  XOR2X1 U29 ( .IN1(A[26]), .IN2(n18), .Q(SUM[26]) );
  XOR2X1 U30 ( .IN1(A[25]), .IN2(n17), .Q(SUM[25]) );
  XOR2X1 U31 ( .IN1(A[24]), .IN2(n16), .Q(SUM[24]) );
  XOR2X1 U32 ( .IN1(A[23]), .IN2(n15), .Q(SUM[23]) );
  XOR2X1 U33 ( .IN1(A[22]), .IN2(n14), .Q(SUM[22]) );
  XOR2X1 U34 ( .IN1(A[21]), .IN2(n13), .Q(SUM[21]) );
  XOR2X1 U35 ( .IN1(A[20]), .IN2(n12), .Q(SUM[20]) );
  XOR2X1 U36 ( .IN1(A[19]), .IN2(n11), .Q(SUM[19]) );
  XOR2X1 U37 ( .IN1(A[18]), .IN2(n10), .Q(SUM[18]) );
  XOR2X1 U38 ( .IN1(A[17]), .IN2(n9), .Q(SUM[17]) );
  XOR2X1 U39 ( .IN1(A[16]), .IN2(n8), .Q(SUM[16]) );
  XOR2X1 U40 ( .IN1(A[15]), .IN2(n7), .Q(SUM[15]) );
  XOR2X1 U41 ( .IN1(A[14]), .IN2(n6), .Q(SUM[14]) );
  XOR2X1 U42 ( .IN1(A[13]), .IN2(n5), .Q(SUM[13]) );
  XOR2X1 U43 ( .IN1(A[12]), .IN2(n4), .Q(SUM[12]) );
  XOR2X1 U44 ( .IN1(A[11]), .IN2(n3), .Q(SUM[11]) );
  XOR2X1 U45 ( .IN1(A[10]), .IN2(carry[10]), .Q(SUM[10]) );
  XOR2X1 U46 ( .IN1(A[2]), .IN2(B[2]), .Q(SUM[2]) );
endmodule


module thumb_DW01_add_2 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [32:1] carry;

  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(n2), .CO(carry[4]), .S(SUM[3]) );
  AND2X1 U1 ( .IN1(A[31]), .IN2(n23), .Q(SUM[32]) );
  AND2X1 U2 ( .IN1(A[2]), .IN2(B[2]), .Q(n2) );
  AND2X1 U3 ( .IN1(A[10]), .IN2(carry[10]), .Q(n3) );
  AND2X1 U4 ( .IN1(A[11]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(A[12]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(A[13]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(A[14]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(A[15]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(A[16]), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(A[17]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(A[18]), .IN2(n10), .Q(n11) );
  AND2X1 U12 ( .IN1(A[19]), .IN2(n11), .Q(n12) );
  AND2X1 U13 ( .IN1(A[20]), .IN2(n12), .Q(n13) );
  AND2X1 U14 ( .IN1(A[21]), .IN2(n13), .Q(n14) );
  AND2X1 U15 ( .IN1(A[22]), .IN2(n14), .Q(n15) );
  AND2X1 U16 ( .IN1(A[23]), .IN2(n15), .Q(n16) );
  AND2X1 U17 ( .IN1(A[24]), .IN2(n16), .Q(n17) );
  AND2X1 U18 ( .IN1(A[25]), .IN2(n17), .Q(n18) );
  AND2X1 U19 ( .IN1(A[26]), .IN2(n18), .Q(n19) );
  AND2X1 U20 ( .IN1(A[27]), .IN2(n19), .Q(n20) );
  AND2X1 U21 ( .IN1(A[28]), .IN2(n20), .Q(n21) );
  AND2X1 U22 ( .IN1(A[29]), .IN2(n21), .Q(n22) );
  AND2X1 U23 ( .IN1(A[30]), .IN2(n22), .Q(n23) );
  XOR2X1 U24 ( .IN1(A[31]), .IN2(n23), .Q(SUM[31]) );
  XOR2X1 U25 ( .IN1(A[30]), .IN2(n22), .Q(SUM[30]) );
  XOR2X1 U26 ( .IN1(A[29]), .IN2(n21), .Q(SUM[29]) );
  XOR2X1 U27 ( .IN1(A[28]), .IN2(n20), .Q(SUM[28]) );
  XOR2X1 U28 ( .IN1(A[27]), .IN2(n19), .Q(SUM[27]) );
  XOR2X1 U29 ( .IN1(A[26]), .IN2(n18), .Q(SUM[26]) );
  XOR2X1 U30 ( .IN1(A[25]), .IN2(n17), .Q(SUM[25]) );
  XOR2X1 U31 ( .IN1(A[24]), .IN2(n16), .Q(SUM[24]) );
  XOR2X1 U32 ( .IN1(A[23]), .IN2(n15), .Q(SUM[23]) );
  XOR2X1 U33 ( .IN1(A[22]), .IN2(n14), .Q(SUM[22]) );
  XOR2X1 U34 ( .IN1(A[21]), .IN2(n13), .Q(SUM[21]) );
  XOR2X1 U35 ( .IN1(A[20]), .IN2(n12), .Q(SUM[20]) );
  XOR2X1 U36 ( .IN1(A[19]), .IN2(n11), .Q(SUM[19]) );
  XOR2X1 U37 ( .IN1(A[18]), .IN2(n10), .Q(SUM[18]) );
  XOR2X1 U38 ( .IN1(A[17]), .IN2(n9), .Q(SUM[17]) );
  XOR2X1 U39 ( .IN1(A[16]), .IN2(n8), .Q(SUM[16]) );
  XOR2X1 U40 ( .IN1(A[15]), .IN2(n7), .Q(SUM[15]) );
  XOR2X1 U41 ( .IN1(A[14]), .IN2(n6), .Q(SUM[14]) );
  XOR2X1 U42 ( .IN1(A[13]), .IN2(n5), .Q(SUM[13]) );
  XOR2X1 U43 ( .IN1(A[12]), .IN2(n4), .Q(SUM[12]) );
  XOR2X1 U44 ( .IN1(A[11]), .IN2(n3), .Q(SUM[11]) );
  XOR2X1 U45 ( .IN1(A[10]), .IN2(carry[10]), .Q(SUM[10]) );
  XOR2X1 U46 ( .IN1(A[2]), .IN2(B[2]), .Q(SUM[2]) );
endmodule


module thumb_DW01_add_3 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [32:1] carry;

  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(SUM[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module thumb_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29;
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  XNOR2X1 U1 ( .IN1(A[31]), .IN2(n29), .Q(SUM[31]) );
  NAND2X1 U2 ( .IN1(A[30]), .IN2(n28), .QN(n29) );
  AND2X1 U3 ( .IN1(A[2]), .IN2(A[1]), .Q(n1) );
  AND2X1 U4 ( .IN1(A[3]), .IN2(n1), .Q(n2) );
  AND2X1 U5 ( .IN1(A[4]), .IN2(n2), .Q(n3) );
  AND2X1 U6 ( .IN1(A[5]), .IN2(n3), .Q(n4) );
  AND2X1 U7 ( .IN1(A[6]), .IN2(n4), .Q(n5) );
  AND2X1 U8 ( .IN1(A[7]), .IN2(n5), .Q(n6) );
  AND2X1 U9 ( .IN1(A[8]), .IN2(n6), .Q(n7) );
  AND2X1 U10 ( .IN1(A[9]), .IN2(n7), .Q(n8) );
  AND2X1 U11 ( .IN1(A[10]), .IN2(n8), .Q(n9) );
  AND2X1 U12 ( .IN1(A[11]), .IN2(n9), .Q(n10) );
  AND2X1 U13 ( .IN1(A[12]), .IN2(n10), .Q(n11) );
  AND2X1 U14 ( .IN1(A[13]), .IN2(n11), .Q(n12) );
  AND2X1 U15 ( .IN1(A[14]), .IN2(n12), .Q(n13) );
  AND2X1 U16 ( .IN1(A[15]), .IN2(n13), .Q(n14) );
  AND2X1 U17 ( .IN1(A[16]), .IN2(n14), .Q(n15) );
  AND2X1 U18 ( .IN1(A[17]), .IN2(n15), .Q(n16) );
  AND2X1 U19 ( .IN1(A[18]), .IN2(n16), .Q(n17) );
  AND2X1 U20 ( .IN1(A[19]), .IN2(n17), .Q(n18) );
  AND2X1 U21 ( .IN1(A[20]), .IN2(n18), .Q(n19) );
  AND2X1 U22 ( .IN1(A[21]), .IN2(n19), .Q(n20) );
  AND2X1 U23 ( .IN1(A[22]), .IN2(n20), .Q(n21) );
  AND2X1 U24 ( .IN1(A[23]), .IN2(n21), .Q(n22) );
  AND2X1 U25 ( .IN1(A[24]), .IN2(n22), .Q(n23) );
  AND2X1 U26 ( .IN1(A[25]), .IN2(n23), .Q(n24) );
  AND2X1 U27 ( .IN1(A[26]), .IN2(n24), .Q(n25) );
  AND2X1 U28 ( .IN1(A[27]), .IN2(n25), .Q(n26) );
  AND2X1 U29 ( .IN1(A[28]), .IN2(n26), .Q(n27) );
  AND2X1 U30 ( .IN1(A[29]), .IN2(n27), .Q(n28) );
  XOR2X1 U31 ( .IN1(A[30]), .IN2(n28), .Q(SUM[30]) );
  XOR2X1 U32 ( .IN1(A[29]), .IN2(n27), .Q(SUM[29]) );
  XOR2X1 U33 ( .IN1(A[28]), .IN2(n26), .Q(SUM[28]) );
  XOR2X1 U34 ( .IN1(A[27]), .IN2(n25), .Q(SUM[27]) );
  XOR2X1 U35 ( .IN1(A[26]), .IN2(n24), .Q(SUM[26]) );
  XOR2X1 U36 ( .IN1(A[25]), .IN2(n23), .Q(SUM[25]) );
  XOR2X1 U37 ( .IN1(A[24]), .IN2(n22), .Q(SUM[24]) );
  XOR2X1 U38 ( .IN1(A[23]), .IN2(n21), .Q(SUM[23]) );
  XOR2X1 U39 ( .IN1(A[22]), .IN2(n20), .Q(SUM[22]) );
  XOR2X1 U40 ( .IN1(A[21]), .IN2(n19), .Q(SUM[21]) );
  XOR2X1 U41 ( .IN1(A[20]), .IN2(n18), .Q(SUM[20]) );
  XOR2X1 U42 ( .IN1(A[19]), .IN2(n17), .Q(SUM[19]) );
  XOR2X1 U43 ( .IN1(A[18]), .IN2(n16), .Q(SUM[18]) );
  XOR2X1 U44 ( .IN1(A[17]), .IN2(n15), .Q(SUM[17]) );
  XOR2X1 U45 ( .IN1(A[16]), .IN2(n14), .Q(SUM[16]) );
  XOR2X1 U46 ( .IN1(A[15]), .IN2(n13), .Q(SUM[15]) );
  XOR2X1 U47 ( .IN1(A[14]), .IN2(n12), .Q(SUM[14]) );
  XOR2X1 U48 ( .IN1(A[13]), .IN2(n11), .Q(SUM[13]) );
  XOR2X1 U49 ( .IN1(A[12]), .IN2(n10), .Q(SUM[12]) );
  XOR2X1 U50 ( .IN1(A[11]), .IN2(n9), .Q(SUM[11]) );
  XOR2X1 U51 ( .IN1(A[10]), .IN2(n8), .Q(SUM[10]) );
  XOR2X1 U52 ( .IN1(A[9]), .IN2(n7), .Q(SUM[9]) );
  XOR2X1 U53 ( .IN1(A[8]), .IN2(n6), .Q(SUM[8]) );
  XOR2X1 U54 ( .IN1(A[7]), .IN2(n5), .Q(SUM[7]) );
  XOR2X1 U55 ( .IN1(A[6]), .IN2(n4), .Q(SUM[6]) );
  XOR2X1 U56 ( .IN1(A[5]), .IN2(n3), .Q(SUM[5]) );
  XOR2X1 U57 ( .IN1(A[4]), .IN2(n2), .Q(SUM[4]) );
  XOR2X1 U58 ( .IN1(A[3]), .IN2(n1), .Q(SUM[3]) );
  XOR2X1 U59 ( .IN1(A[2]), .IN2(A[1]), .Q(SUM[2]) );
  INVX0 U60 ( .INP(A[1]), .ZN(SUM[1]) );
endmodule


module thumb_DW_leftsh_2 ( A, SH, B );
  input [32:0] A;
  input [4:0] SH;
  output [32:0] B;
  wire   n1, n17, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163;

  MUX21X1 U1 ( .IN1(n57), .IN2(n41), .S(SH[4]), .Q(B[32]) );
  MUX21X1 U2 ( .IN1(n56), .IN2(n40), .S(SH[4]), .Q(B[31]) );
  MUX21X1 U3 ( .IN1(n55), .IN2(n39), .S(SH[4]), .Q(B[30]) );
  MUX21X1 U4 ( .IN1(n54), .IN2(n38), .S(SH[4]), .Q(B[29]) );
  MUX21X1 U5 ( .IN1(n53), .IN2(n37), .S(SH[4]), .Q(B[28]) );
  MUX21X1 U6 ( .IN1(n52), .IN2(n36), .S(SH[4]), .Q(B[27]) );
  MUX21X1 U7 ( .IN1(n51), .IN2(n35), .S(SH[4]), .Q(B[26]) );
  MUX21X1 U8 ( .IN1(n50), .IN2(n34), .S(SH[4]), .Q(B[25]) );
  MUX21X1 U9 ( .IN1(n49), .IN2(n33), .S(SH[4]), .Q(B[24]) );
  MUX21X1 U10 ( .IN1(n48), .IN2(n32), .S(SH[4]), .Q(B[23]) );
  MUX21X1 U11 ( .IN1(n47), .IN2(n31), .S(SH[4]), .Q(B[22]) );
  MUX21X1 U12 ( .IN1(n46), .IN2(n30), .S(SH[4]), .Q(B[21]) );
  MUX21X1 U13 ( .IN1(n45), .IN2(n29), .S(SH[4]), .Q(B[20]) );
  MUX21X1 U14 ( .IN1(n44), .IN2(n28), .S(SH[4]), .Q(B[19]) );
  MUX21X1 U15 ( .IN1(n43), .IN2(n27), .S(SH[4]), .Q(B[18]) );
  MUX21X1 U16 ( .IN1(n42), .IN2(n26), .S(SH[4]), .Q(B[17]) );
  MUX21X1 U17 ( .IN1(n41), .IN2(n25), .S(SH[4]), .Q(B[16]) );
  MUX21X1 U50 ( .IN1(n94), .IN2(n86), .S(SH[3]), .Q(n57) );
  MUX21X1 U51 ( .IN1(n93), .IN2(n85), .S(SH[3]), .Q(n56) );
  MUX21X1 U52 ( .IN1(n92), .IN2(n84), .S(SH[3]), .Q(n55) );
  MUX21X1 U53 ( .IN1(n91), .IN2(n83), .S(SH[3]), .Q(n54) );
  MUX21X1 U54 ( .IN1(n90), .IN2(n82), .S(SH[3]), .Q(n53) );
  MUX21X1 U55 ( .IN1(n89), .IN2(n81), .S(SH[3]), .Q(n52) );
  MUX21X1 U56 ( .IN1(n88), .IN2(n80), .S(SH[3]), .Q(n51) );
  MUX21X1 U57 ( .IN1(n87), .IN2(n79), .S(SH[3]), .Q(n50) );
  MUX21X1 U58 ( .IN1(n86), .IN2(n78), .S(SH[3]), .Q(n49) );
  MUX21X1 U59 ( .IN1(n85), .IN2(n77), .S(SH[3]), .Q(n48) );
  MUX21X1 U60 ( .IN1(n84), .IN2(n76), .S(SH[3]), .Q(n47) );
  MUX21X1 U61 ( .IN1(n83), .IN2(n75), .S(SH[3]), .Q(n46) );
  MUX21X1 U62 ( .IN1(n82), .IN2(n74), .S(SH[3]), .Q(n45) );
  MUX21X1 U63 ( .IN1(n81), .IN2(n73), .S(SH[3]), .Q(n44) );
  MUX21X1 U64 ( .IN1(n80), .IN2(n72), .S(SH[3]), .Q(n43) );
  MUX21X1 U65 ( .IN1(n79), .IN2(n71), .S(SH[3]), .Q(n42) );
  MUX21X1 U66 ( .IN1(n78), .IN2(n70), .S(SH[3]), .Q(n41) );
  MUX21X1 U67 ( .IN1(n77), .IN2(n69), .S(SH[3]), .Q(n40) );
  MUX21X1 U68 ( .IN1(n76), .IN2(n68), .S(SH[3]), .Q(n39) );
  MUX21X1 U69 ( .IN1(n75), .IN2(n67), .S(SH[3]), .Q(n38) );
  MUX21X1 U70 ( .IN1(n74), .IN2(n66), .S(SH[3]), .Q(n37) );
  MUX21X1 U71 ( .IN1(n73), .IN2(n65), .S(SH[3]), .Q(n36) );
  MUX21X1 U72 ( .IN1(n72), .IN2(n64), .S(SH[3]), .Q(n35) );
  MUX21X1 U73 ( .IN1(n71), .IN2(n63), .S(SH[3]), .Q(n34) );
  MUX21X1 U74 ( .IN1(n70), .IN2(n62), .S(SH[3]), .Q(n33) );
  MUX21X1 U91 ( .IN1(n129), .IN2(n125), .S(SH[2]), .Q(n94) );
  MUX21X1 U92 ( .IN1(n128), .IN2(n124), .S(SH[2]), .Q(n93) );
  MUX21X1 U93 ( .IN1(n127), .IN2(n123), .S(SH[2]), .Q(n92) );
  MUX21X1 U94 ( .IN1(n126), .IN2(n122), .S(SH[2]), .Q(n91) );
  MUX21X1 U95 ( .IN1(n125), .IN2(n121), .S(SH[2]), .Q(n90) );
  MUX21X1 U96 ( .IN1(n124), .IN2(n120), .S(SH[2]), .Q(n89) );
  MUX21X1 U97 ( .IN1(n123), .IN2(n119), .S(SH[2]), .Q(n88) );
  MUX21X1 U98 ( .IN1(n122), .IN2(n118), .S(SH[2]), .Q(n87) );
  MUX21X1 U99 ( .IN1(n121), .IN2(n117), .S(SH[2]), .Q(n86) );
  MUX21X1 U100 ( .IN1(n120), .IN2(n116), .S(SH[2]), .Q(n85) );
  MUX21X1 U101 ( .IN1(n119), .IN2(n115), .S(SH[2]), .Q(n84) );
  MUX21X1 U102 ( .IN1(n118), .IN2(n114), .S(SH[2]), .Q(n83) );
  MUX21X1 U103 ( .IN1(n117), .IN2(n113), .S(SH[2]), .Q(n82) );
  MUX21X1 U104 ( .IN1(n116), .IN2(n112), .S(SH[2]), .Q(n81) );
  MUX21X1 U105 ( .IN1(n115), .IN2(n111), .S(SH[2]), .Q(n80) );
  MUX21X1 U106 ( .IN1(n114), .IN2(n110), .S(SH[2]), .Q(n79) );
  MUX21X1 U107 ( .IN1(n113), .IN2(n109), .S(SH[2]), .Q(n78) );
  MUX21X1 U108 ( .IN1(n112), .IN2(n108), .S(SH[2]), .Q(n77) );
  MUX21X1 U109 ( .IN1(n111), .IN2(n107), .S(SH[2]), .Q(n76) );
  MUX21X1 U110 ( .IN1(n110), .IN2(n106), .S(SH[2]), .Q(n75) );
  MUX21X1 U111 ( .IN1(n109), .IN2(n105), .S(SH[2]), .Q(n74) );
  MUX21X1 U112 ( .IN1(n108), .IN2(n104), .S(SH[2]), .Q(n73) );
  MUX21X1 U113 ( .IN1(n107), .IN2(n103), .S(SH[2]), .Q(n72) );
  MUX21X1 U114 ( .IN1(n106), .IN2(n102), .S(SH[2]), .Q(n71) );
  MUX21X1 U115 ( .IN1(n105), .IN2(n101), .S(SH[2]), .Q(n70) );
  MUX21X1 U116 ( .IN1(n104), .IN2(n100), .S(SH[2]), .Q(n69) );
  MUX21X1 U117 ( .IN1(n103), .IN2(n99), .S(SH[2]), .Q(n68) );
  MUX21X1 U118 ( .IN1(n102), .IN2(n98), .S(SH[2]), .Q(n67) );
  MUX21X1 U119 ( .IN1(n101), .IN2(n97), .S(SH[2]), .Q(n66) );
  MUX21X1 U128 ( .IN1(n163), .IN2(n161), .S(SH[1]), .Q(n129) );
  MUX21X1 U129 ( .IN1(n162), .IN2(n160), .S(SH[1]), .Q(n128) );
  MUX21X1 U130 ( .IN1(n161), .IN2(n159), .S(SH[1]), .Q(n127) );
  MUX21X1 U131 ( .IN1(n160), .IN2(n158), .S(SH[1]), .Q(n126) );
  MUX21X1 U132 ( .IN1(n159), .IN2(n157), .S(SH[1]), .Q(n125) );
  MUX21X1 U133 ( .IN1(n158), .IN2(n156), .S(SH[1]), .Q(n124) );
  MUX21X1 U134 ( .IN1(n157), .IN2(n155), .S(SH[1]), .Q(n123) );
  MUX21X1 U135 ( .IN1(n156), .IN2(n154), .S(SH[1]), .Q(n122) );
  MUX21X1 U136 ( .IN1(n155), .IN2(n153), .S(SH[1]), .Q(n121) );
  MUX21X1 U137 ( .IN1(n154), .IN2(n152), .S(SH[1]), .Q(n120) );
  MUX21X1 U138 ( .IN1(n153), .IN2(n151), .S(SH[1]), .Q(n119) );
  MUX21X1 U139 ( .IN1(n152), .IN2(n150), .S(SH[1]), .Q(n118) );
  MUX21X1 U140 ( .IN1(n151), .IN2(n149), .S(SH[1]), .Q(n117) );
  MUX21X1 U141 ( .IN1(n150), .IN2(n148), .S(SH[1]), .Q(n116) );
  MUX21X1 U142 ( .IN1(n149), .IN2(n147), .S(SH[1]), .Q(n115) );
  MUX21X1 U143 ( .IN1(n148), .IN2(n146), .S(SH[1]), .Q(n114) );
  MUX21X1 U144 ( .IN1(n147), .IN2(n145), .S(SH[1]), .Q(n113) );
  MUX21X1 U145 ( .IN1(n146), .IN2(n144), .S(SH[1]), .Q(n112) );
  MUX21X1 U146 ( .IN1(n145), .IN2(n143), .S(SH[1]), .Q(n111) );
  MUX21X1 U147 ( .IN1(n144), .IN2(n142), .S(SH[1]), .Q(n110) );
  MUX21X1 U148 ( .IN1(n143), .IN2(n141), .S(SH[1]), .Q(n109) );
  MUX21X1 U149 ( .IN1(n142), .IN2(n140), .S(SH[1]), .Q(n108) );
  MUX21X1 U150 ( .IN1(n141), .IN2(n139), .S(SH[1]), .Q(n107) );
  MUX21X1 U151 ( .IN1(n140), .IN2(n138), .S(SH[1]), .Q(n106) );
  MUX21X1 U152 ( .IN1(n139), .IN2(n137), .S(SH[1]), .Q(n105) );
  MUX21X1 U153 ( .IN1(n138), .IN2(n136), .S(SH[1]), .Q(n104) );
  MUX21X1 U154 ( .IN1(n137), .IN2(n135), .S(SH[1]), .Q(n103) );
  MUX21X1 U155 ( .IN1(n136), .IN2(n134), .S(SH[1]), .Q(n102) );
  MUX21X1 U156 ( .IN1(n135), .IN2(n133), .S(SH[1]), .Q(n101) );
  MUX21X1 U157 ( .IN1(n134), .IN2(n132), .S(SH[1]), .Q(n100) );
  MUX21X1 U158 ( .IN1(n133), .IN2(n131), .S(SH[1]), .Q(n99) );
  AND2X1 U163 ( .IN1(SH[0]), .IN2(A[31]), .Q(n163) );
  MUX21X1 U164 ( .IN1(A[31]), .IN2(A[30]), .S(SH[0]), .Q(n162) );
  MUX21X1 U165 ( .IN1(A[30]), .IN2(A[29]), .S(SH[0]), .Q(n161) );
  MUX21X1 U166 ( .IN1(A[29]), .IN2(A[28]), .S(SH[0]), .Q(n160) );
  MUX21X1 U167 ( .IN1(A[28]), .IN2(A[27]), .S(SH[0]), .Q(n159) );
  MUX21X1 U168 ( .IN1(A[27]), .IN2(A[26]), .S(SH[0]), .Q(n158) );
  MUX21X1 U169 ( .IN1(A[26]), .IN2(A[25]), .S(SH[0]), .Q(n157) );
  MUX21X1 U170 ( .IN1(A[25]), .IN2(A[24]), .S(SH[0]), .Q(n156) );
  MUX21X1 U171 ( .IN1(A[24]), .IN2(A[23]), .S(SH[0]), .Q(n155) );
  MUX21X1 U172 ( .IN1(A[23]), .IN2(A[22]), .S(SH[0]), .Q(n154) );
  MUX21X1 U173 ( .IN1(A[22]), .IN2(A[21]), .S(SH[0]), .Q(n153) );
  MUX21X1 U174 ( .IN1(A[21]), .IN2(A[20]), .S(SH[0]), .Q(n152) );
  MUX21X1 U175 ( .IN1(A[20]), .IN2(A[19]), .S(SH[0]), .Q(n151) );
  MUX21X1 U176 ( .IN1(A[19]), .IN2(A[18]), .S(SH[0]), .Q(n150) );
  MUX21X1 U177 ( .IN1(A[18]), .IN2(A[17]), .S(SH[0]), .Q(n149) );
  MUX21X1 U178 ( .IN1(A[17]), .IN2(A[16]), .S(SH[0]), .Q(n148) );
  MUX21X1 U179 ( .IN1(A[16]), .IN2(A[15]), .S(SH[0]), .Q(n147) );
  MUX21X1 U180 ( .IN1(A[15]), .IN2(A[14]), .S(SH[0]), .Q(n146) );
  MUX21X1 U181 ( .IN1(A[14]), .IN2(A[13]), .S(SH[0]), .Q(n145) );
  MUX21X1 U182 ( .IN1(A[13]), .IN2(A[12]), .S(SH[0]), .Q(n144) );
  MUX21X1 U183 ( .IN1(A[12]), .IN2(A[11]), .S(SH[0]), .Q(n143) );
  MUX21X1 U184 ( .IN1(A[11]), .IN2(A[10]), .S(SH[0]), .Q(n142) );
  MUX21X1 U185 ( .IN1(A[10]), .IN2(A[9]), .S(SH[0]), .Q(n141) );
  MUX21X1 U186 ( .IN1(A[9]), .IN2(A[8]), .S(SH[0]), .Q(n140) );
  MUX21X1 U187 ( .IN1(A[8]), .IN2(A[7]), .S(SH[0]), .Q(n139) );
  MUX21X1 U188 ( .IN1(A[7]), .IN2(A[6]), .S(SH[0]), .Q(n138) );
  MUX21X1 U189 ( .IN1(A[6]), .IN2(A[5]), .S(SH[0]), .Q(n137) );
  MUX21X1 U190 ( .IN1(A[5]), .IN2(A[4]), .S(SH[0]), .Q(n136) );
  MUX21X1 U191 ( .IN1(A[4]), .IN2(A[3]), .S(SH[0]), .Q(n135) );
  MUX21X1 U192 ( .IN1(A[3]), .IN2(A[2]), .S(SH[0]), .Q(n134) );
  MUX21X1 U193 ( .IN1(A[2]), .IN2(A[1]), .S(SH[0]), .Q(n133) );
  MUX21X1 U194 ( .IN1(A[1]), .IN2(A[0]), .S(SH[0]), .Q(n132) );
  AND2X1 U200 ( .IN1(n40), .IN2(n1), .Q(B[15]) );
  AND2X1 U201 ( .IN1(n39), .IN2(n1), .Q(B[14]) );
  AND2X1 U202 ( .IN1(n38), .IN2(n1), .Q(B[13]) );
  AND2X1 U203 ( .IN1(n37), .IN2(n1), .Q(B[12]) );
  AND2X1 U204 ( .IN1(n36), .IN2(n1), .Q(B[11]) );
  AND2X1 U205 ( .IN1(n35), .IN2(n1), .Q(B[10]) );
  AND2X1 U206 ( .IN1(n34), .IN2(n1), .Q(B[9]) );
  AND2X1 U207 ( .IN1(n33), .IN2(n1), .Q(B[8]) );
  AND2X1 U208 ( .IN1(n32), .IN2(n1), .Q(B[7]) );
  AND2X1 U209 ( .IN1(n31), .IN2(n1), .Q(B[6]) );
  AND2X1 U210 ( .IN1(n30), .IN2(n1), .Q(B[5]) );
  AND2X1 U211 ( .IN1(n29), .IN2(n1), .Q(B[4]) );
  AND2X1 U212 ( .IN1(n28), .IN2(n1), .Q(B[3]) );
  AND2X1 U213 ( .IN1(n27), .IN2(n1), .Q(B[2]) );
  AND2X1 U214 ( .IN1(n26), .IN2(n1), .Q(B[1]) );
  AND2X1 U215 ( .IN1(n25), .IN2(n1), .Q(B[0]) );
  AND2X1 U216 ( .IN1(n69), .IN2(n17), .Q(n32) );
  AND2X1 U217 ( .IN1(n68), .IN2(n17), .Q(n31) );
  AND2X1 U218 ( .IN1(n67), .IN2(n17), .Q(n30) );
  AND2X1 U219 ( .IN1(n66), .IN2(n17), .Q(n29) );
  AND2X1 U220 ( .IN1(n65), .IN2(n17), .Q(n28) );
  AND2X1 U221 ( .IN1(n64), .IN2(n17), .Q(n27) );
  AND2X1 U222 ( .IN1(n63), .IN2(n17), .Q(n26) );
  AND2X1 U223 ( .IN1(n62), .IN2(n17), .Q(n25) );
  AND2X1 U224 ( .IN1(n100), .IN2(n58), .Q(n65) );
  AND2X1 U225 ( .IN1(n99), .IN2(n58), .Q(n64) );
  AND2X1 U226 ( .IN1(n98), .IN2(n58), .Q(n63) );
  AND2X1 U227 ( .IN1(n97), .IN2(n58), .Q(n62) );
  AND2X1 U228 ( .IN1(n132), .IN2(n95), .Q(n98) );
  AND2X1 U229 ( .IN1(n131), .IN2(n95), .Q(n97) );
  INVX0 U230 ( .INP(SH[4]), .ZN(n1) );
  INVX0 U231 ( .INP(SH[3]), .ZN(n17) );
  INVX0 U232 ( .INP(SH[2]), .ZN(n58) );
  INVX0 U233 ( .INP(SH[1]), .ZN(n95) );
  AND2X1 U234 ( .IN1(A[0]), .IN2(n130), .Q(n131) );
  INVX0 U235 ( .INP(SH[0]), .ZN(n130) );
endmodule


module thumb_DW_rightsh_2 ( A, DATA_TC, SH, B );
  input [32:0] A;
  input [4:0] SH;
  output [32:0] B;
  input DATA_TC;
  wire   n1, n17, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163;

  MUX21X1 U33 ( .IN1(n41), .IN2(n57), .S(SH[4]), .Q(B[16]) );
  MUX21X1 U34 ( .IN1(n40), .IN2(n56), .S(SH[4]), .Q(B[15]) );
  MUX21X1 U35 ( .IN1(n39), .IN2(n55), .S(SH[4]), .Q(B[14]) );
  MUX21X1 U36 ( .IN1(n38), .IN2(n54), .S(SH[4]), .Q(B[13]) );
  MUX21X1 U37 ( .IN1(n37), .IN2(n53), .S(SH[4]), .Q(B[12]) );
  MUX21X1 U38 ( .IN1(n36), .IN2(n52), .S(SH[4]), .Q(B[11]) );
  MUX21X1 U39 ( .IN1(n35), .IN2(n51), .S(SH[4]), .Q(B[10]) );
  MUX21X1 U40 ( .IN1(n34), .IN2(n50), .S(SH[4]), .Q(B[9]) );
  MUX21X1 U41 ( .IN1(n33), .IN2(n49), .S(SH[4]), .Q(B[8]) );
  MUX21X1 U42 ( .IN1(n32), .IN2(n48), .S(SH[4]), .Q(B[7]) );
  MUX21X1 U43 ( .IN1(n31), .IN2(n47), .S(SH[4]), .Q(B[6]) );
  MUX21X1 U44 ( .IN1(n30), .IN2(n46), .S(SH[4]), .Q(B[5]) );
  MUX21X1 U45 ( .IN1(n29), .IN2(n45), .S(SH[4]), .Q(B[4]) );
  MUX21X1 U46 ( .IN1(n28), .IN2(n44), .S(SH[4]), .Q(B[3]) );
  MUX21X1 U47 ( .IN1(n27), .IN2(n43), .S(SH[4]), .Q(B[2]) );
  MUX21X1 U48 ( .IN1(n26), .IN2(n42), .S(SH[4]), .Q(B[1]) );
  MUX21X1 U49 ( .IN1(n25), .IN2(n41), .S(SH[4]), .Q(B[0]) );
  MUX21X1 U66 ( .IN1(n86), .IN2(n94), .S(SH[3]), .Q(n49) );
  MUX21X1 U67 ( .IN1(n85), .IN2(n93), .S(SH[3]), .Q(n48) );
  MUX21X1 U68 ( .IN1(n84), .IN2(n92), .S(SH[3]), .Q(n47) );
  MUX21X1 U69 ( .IN1(n83), .IN2(n91), .S(SH[3]), .Q(n46) );
  MUX21X1 U70 ( .IN1(n82), .IN2(n90), .S(SH[3]), .Q(n45) );
  MUX21X1 U71 ( .IN1(n81), .IN2(n89), .S(SH[3]), .Q(n44) );
  MUX21X1 U72 ( .IN1(n80), .IN2(n88), .S(SH[3]), .Q(n43) );
  MUX21X1 U73 ( .IN1(n79), .IN2(n87), .S(SH[3]), .Q(n42) );
  MUX21X1 U74 ( .IN1(n78), .IN2(n86), .S(SH[3]), .Q(n41) );
  MUX21X1 U75 ( .IN1(n77), .IN2(n85), .S(SH[3]), .Q(n40) );
  MUX21X1 U76 ( .IN1(n76), .IN2(n84), .S(SH[3]), .Q(n39) );
  MUX21X1 U77 ( .IN1(n75), .IN2(n83), .S(SH[3]), .Q(n38) );
  MUX21X1 U78 ( .IN1(n74), .IN2(n82), .S(SH[3]), .Q(n37) );
  MUX21X1 U79 ( .IN1(n73), .IN2(n81), .S(SH[3]), .Q(n36) );
  MUX21X1 U80 ( .IN1(n72), .IN2(n80), .S(SH[3]), .Q(n35) );
  MUX21X1 U81 ( .IN1(n71), .IN2(n79), .S(SH[3]), .Q(n34) );
  MUX21X1 U82 ( .IN1(n70), .IN2(n78), .S(SH[3]), .Q(n33) );
  MUX21X1 U83 ( .IN1(n69), .IN2(n77), .S(SH[3]), .Q(n32) );
  MUX21X1 U84 ( .IN1(n68), .IN2(n76), .S(SH[3]), .Q(n31) );
  MUX21X1 U85 ( .IN1(n67), .IN2(n75), .S(SH[3]), .Q(n30) );
  MUX21X1 U86 ( .IN1(n66), .IN2(n74), .S(SH[3]), .Q(n29) );
  MUX21X1 U87 ( .IN1(n65), .IN2(n73), .S(SH[3]), .Q(n28) );
  MUX21X1 U88 ( .IN1(n64), .IN2(n72), .S(SH[3]), .Q(n27) );
  MUX21X1 U89 ( .IN1(n63), .IN2(n71), .S(SH[3]), .Q(n26) );
  MUX21X1 U90 ( .IN1(n62), .IN2(n70), .S(SH[3]), .Q(n25) );
  MUX21X1 U99 ( .IN1(n125), .IN2(n129), .S(SH[2]), .Q(n90) );
  MUX21X1 U100 ( .IN1(n124), .IN2(n128), .S(SH[2]), .Q(n89) );
  MUX21X1 U101 ( .IN1(n123), .IN2(n127), .S(SH[2]), .Q(n88) );
  MUX21X1 U102 ( .IN1(n122), .IN2(n126), .S(SH[2]), .Q(n87) );
  MUX21X1 U103 ( .IN1(n121), .IN2(n125), .S(SH[2]), .Q(n86) );
  MUX21X1 U104 ( .IN1(n120), .IN2(n124), .S(SH[2]), .Q(n85) );
  MUX21X1 U105 ( .IN1(n119), .IN2(n123), .S(SH[2]), .Q(n84) );
  MUX21X1 U106 ( .IN1(n118), .IN2(n122), .S(SH[2]), .Q(n83) );
  MUX21X1 U107 ( .IN1(n117), .IN2(n121), .S(SH[2]), .Q(n82) );
  MUX21X1 U108 ( .IN1(n116), .IN2(n120), .S(SH[2]), .Q(n81) );
  MUX21X1 U109 ( .IN1(n115), .IN2(n119), .S(SH[2]), .Q(n80) );
  MUX21X1 U110 ( .IN1(n114), .IN2(n118), .S(SH[2]), .Q(n79) );
  MUX21X1 U111 ( .IN1(n113), .IN2(n117), .S(SH[2]), .Q(n78) );
  MUX21X1 U112 ( .IN1(n112), .IN2(n116), .S(SH[2]), .Q(n77) );
  MUX21X1 U113 ( .IN1(n111), .IN2(n115), .S(SH[2]), .Q(n76) );
  MUX21X1 U114 ( .IN1(n110), .IN2(n114), .S(SH[2]), .Q(n75) );
  MUX21X1 U115 ( .IN1(n109), .IN2(n113), .S(SH[2]), .Q(n74) );
  MUX21X1 U116 ( .IN1(n108), .IN2(n112), .S(SH[2]), .Q(n73) );
  MUX21X1 U117 ( .IN1(n107), .IN2(n111), .S(SH[2]), .Q(n72) );
  MUX21X1 U118 ( .IN1(n106), .IN2(n110), .S(SH[2]), .Q(n71) );
  MUX21X1 U119 ( .IN1(n105), .IN2(n109), .S(SH[2]), .Q(n70) );
  MUX21X1 U120 ( .IN1(n104), .IN2(n108), .S(SH[2]), .Q(n69) );
  MUX21X1 U121 ( .IN1(n103), .IN2(n107), .S(SH[2]), .Q(n68) );
  MUX21X1 U122 ( .IN1(n102), .IN2(n106), .S(SH[2]), .Q(n67) );
  MUX21X1 U123 ( .IN1(n101), .IN2(n105), .S(SH[2]), .Q(n66) );
  MUX21X1 U124 ( .IN1(n100), .IN2(n104), .S(SH[2]), .Q(n65) );
  MUX21X1 U125 ( .IN1(n99), .IN2(n103), .S(SH[2]), .Q(n64) );
  MUX21X1 U126 ( .IN1(n98), .IN2(n102), .S(SH[2]), .Q(n63) );
  MUX21X1 U127 ( .IN1(n97), .IN2(n101), .S(SH[2]), .Q(n62) );
  MUX21X1 U132 ( .IN1(n161), .IN2(n163), .S(SH[1]), .Q(n127) );
  MUX21X1 U133 ( .IN1(n160), .IN2(n162), .S(SH[1]), .Q(n126) );
  MUX21X1 U134 ( .IN1(n159), .IN2(n161), .S(SH[1]), .Q(n125) );
  MUX21X1 U135 ( .IN1(n158), .IN2(n160), .S(SH[1]), .Q(n124) );
  MUX21X1 U136 ( .IN1(n157), .IN2(n159), .S(SH[1]), .Q(n123) );
  MUX21X1 U137 ( .IN1(n156), .IN2(n158), .S(SH[1]), .Q(n122) );
  MUX21X1 U138 ( .IN1(n155), .IN2(n157), .S(SH[1]), .Q(n121) );
  MUX21X1 U139 ( .IN1(n154), .IN2(n156), .S(SH[1]), .Q(n120) );
  MUX21X1 U140 ( .IN1(n153), .IN2(n155), .S(SH[1]), .Q(n119) );
  MUX21X1 U141 ( .IN1(n152), .IN2(n154), .S(SH[1]), .Q(n118) );
  MUX21X1 U142 ( .IN1(n151), .IN2(n153), .S(SH[1]), .Q(n117) );
  MUX21X1 U143 ( .IN1(n150), .IN2(n152), .S(SH[1]), .Q(n116) );
  MUX21X1 U144 ( .IN1(n149), .IN2(n151), .S(SH[1]), .Q(n115) );
  MUX21X1 U145 ( .IN1(n148), .IN2(n150), .S(SH[1]), .Q(n114) );
  MUX21X1 U146 ( .IN1(n147), .IN2(n149), .S(SH[1]), .Q(n113) );
  MUX21X1 U147 ( .IN1(n146), .IN2(n148), .S(SH[1]), .Q(n112) );
  MUX21X1 U148 ( .IN1(n145), .IN2(n147), .S(SH[1]), .Q(n111) );
  MUX21X1 U149 ( .IN1(n144), .IN2(n146), .S(SH[1]), .Q(n110) );
  MUX21X1 U150 ( .IN1(n143), .IN2(n145), .S(SH[1]), .Q(n109) );
  MUX21X1 U151 ( .IN1(n142), .IN2(n144), .S(SH[1]), .Q(n108) );
  MUX21X1 U152 ( .IN1(n141), .IN2(n143), .S(SH[1]), .Q(n107) );
  MUX21X1 U153 ( .IN1(n140), .IN2(n142), .S(SH[1]), .Q(n106) );
  MUX21X1 U154 ( .IN1(n139), .IN2(n141), .S(SH[1]), .Q(n105) );
  MUX21X1 U155 ( .IN1(n138), .IN2(n140), .S(SH[1]), .Q(n104) );
  MUX21X1 U156 ( .IN1(n137), .IN2(n139), .S(SH[1]), .Q(n103) );
  MUX21X1 U157 ( .IN1(n136), .IN2(n138), .S(SH[1]), .Q(n102) );
  MUX21X1 U158 ( .IN1(n135), .IN2(n137), .S(SH[1]), .Q(n101) );
  MUX21X1 U159 ( .IN1(n134), .IN2(n136), .S(SH[1]), .Q(n100) );
  MUX21X1 U160 ( .IN1(n133), .IN2(n135), .S(SH[1]), .Q(n99) );
  MUX21X1 U161 ( .IN1(n132), .IN2(n134), .S(SH[1]), .Q(n98) );
  MUX21X1 U162 ( .IN1(n131), .IN2(n133), .S(SH[1]), .Q(n97) );
  MUX21X1 U165 ( .IN1(A[31]), .IN2(A[32]), .S(SH[0]), .Q(n162) );
  MUX21X1 U166 ( .IN1(A[30]), .IN2(A[31]), .S(SH[0]), .Q(n161) );
  MUX21X1 U167 ( .IN1(A[29]), .IN2(A[30]), .S(SH[0]), .Q(n160) );
  MUX21X1 U168 ( .IN1(A[28]), .IN2(A[29]), .S(SH[0]), .Q(n159) );
  MUX21X1 U169 ( .IN1(A[27]), .IN2(A[28]), .S(SH[0]), .Q(n158) );
  MUX21X1 U170 ( .IN1(A[26]), .IN2(A[27]), .S(SH[0]), .Q(n157) );
  MUX21X1 U171 ( .IN1(A[25]), .IN2(A[26]), .S(SH[0]), .Q(n156) );
  MUX21X1 U172 ( .IN1(A[24]), .IN2(A[25]), .S(SH[0]), .Q(n155) );
  MUX21X1 U173 ( .IN1(A[23]), .IN2(A[24]), .S(SH[0]), .Q(n154) );
  MUX21X1 U174 ( .IN1(A[22]), .IN2(A[23]), .S(SH[0]), .Q(n153) );
  MUX21X1 U175 ( .IN1(A[21]), .IN2(A[22]), .S(SH[0]), .Q(n152) );
  MUX21X1 U176 ( .IN1(A[20]), .IN2(A[21]), .S(SH[0]), .Q(n151) );
  MUX21X1 U177 ( .IN1(A[19]), .IN2(A[20]), .S(SH[0]), .Q(n150) );
  MUX21X1 U178 ( .IN1(A[18]), .IN2(A[19]), .S(SH[0]), .Q(n149) );
  MUX21X1 U179 ( .IN1(A[17]), .IN2(A[18]), .S(SH[0]), .Q(n148) );
  MUX21X1 U180 ( .IN1(A[16]), .IN2(A[17]), .S(SH[0]), .Q(n147) );
  MUX21X1 U181 ( .IN1(A[15]), .IN2(A[16]), .S(SH[0]), .Q(n146) );
  MUX21X1 U182 ( .IN1(A[14]), .IN2(A[15]), .S(SH[0]), .Q(n145) );
  MUX21X1 U183 ( .IN1(A[13]), .IN2(A[14]), .S(SH[0]), .Q(n144) );
  MUX21X1 U184 ( .IN1(A[12]), .IN2(A[13]), .S(SH[0]), .Q(n143) );
  MUX21X1 U185 ( .IN1(A[11]), .IN2(A[12]), .S(SH[0]), .Q(n142) );
  MUX21X1 U186 ( .IN1(A[10]), .IN2(A[11]), .S(SH[0]), .Q(n141) );
  MUX21X1 U187 ( .IN1(A[9]), .IN2(A[10]), .S(SH[0]), .Q(n140) );
  MUX21X1 U188 ( .IN1(A[8]), .IN2(A[9]), .S(SH[0]), .Q(n139) );
  MUX21X1 U189 ( .IN1(A[7]), .IN2(A[8]), .S(SH[0]), .Q(n138) );
  MUX21X1 U190 ( .IN1(A[6]), .IN2(A[7]), .S(SH[0]), .Q(n137) );
  MUX21X1 U191 ( .IN1(A[5]), .IN2(A[6]), .S(SH[0]), .Q(n136) );
  MUX21X1 U192 ( .IN1(A[4]), .IN2(A[5]), .S(SH[0]), .Q(n135) );
  MUX21X1 U193 ( .IN1(A[3]), .IN2(A[4]), .S(SH[0]), .Q(n134) );
  MUX21X1 U194 ( .IN1(A[2]), .IN2(A[3]), .S(SH[0]), .Q(n133) );
  MUX21X1 U195 ( .IN1(A[1]), .IN2(A[2]), .S(SH[0]), .Q(n132) );
  AND2X1 U196 ( .IN1(SH[0]), .IN2(A[1]), .Q(n131) );
  AND2X1 U200 ( .IN1(n53), .IN2(n1), .Q(B[28]) );
  AND2X1 U201 ( .IN1(n52), .IN2(n1), .Q(B[27]) );
  AND2X1 U202 ( .IN1(n93), .IN2(n17), .Q(n56) );
  AND2X1 U203 ( .IN1(n92), .IN2(n17), .Q(n55) );
  AND2X1 U204 ( .IN1(n91), .IN2(n17), .Q(n54) );
  AND2X1 U205 ( .IN1(n94), .IN2(n17), .Q(n57) );
  AND2X1 U206 ( .IN1(n90), .IN2(n17), .Q(n53) );
  AND2X1 U207 ( .IN1(n89), .IN2(n17), .Q(n52) );
  AND2X1 U208 ( .IN1(n88), .IN2(n17), .Q(n51) );
  AND2X1 U209 ( .IN1(n87), .IN2(n17), .Q(n50) );
  AND2X1 U210 ( .IN1(n128), .IN2(n58), .Q(n93) );
  AND2X1 U211 ( .IN1(n127), .IN2(n58), .Q(n92) );
  AND2X1 U212 ( .IN1(n126), .IN2(n58), .Q(n91) );
  AND2X1 U213 ( .IN1(n129), .IN2(n58), .Q(n94) );
  AND2X1 U214 ( .IN1(n162), .IN2(n95), .Q(n128) );
  AND2X1 U215 ( .IN1(n163), .IN2(n95), .Q(n129) );
  AND2X1 U216 ( .IN1(n57), .IN2(n1), .Q(B[32]) );
  AND2X1 U217 ( .IN1(n51), .IN2(n1), .Q(B[26]) );
  AND2X1 U218 ( .IN1(n50), .IN2(n1), .Q(B[25]) );
  AND2X1 U219 ( .IN1(n49), .IN2(n1), .Q(B[24]) );
  AND2X1 U220 ( .IN1(n48), .IN2(n1), .Q(B[23]) );
  AND2X1 U221 ( .IN1(n47), .IN2(n1), .Q(B[22]) );
  AND2X1 U222 ( .IN1(n46), .IN2(n1), .Q(B[21]) );
  AND2X1 U223 ( .IN1(n45), .IN2(n1), .Q(B[20]) );
  AND2X1 U224 ( .IN1(n44), .IN2(n1), .Q(B[19]) );
  AND2X1 U225 ( .IN1(n43), .IN2(n1), .Q(B[18]) );
  AND2X1 U226 ( .IN1(n42), .IN2(n1), .Q(B[17]) );
  AND2X1 U227 ( .IN1(n54), .IN2(n1), .Q(B[29]) );
  INVX0 U228 ( .INP(SH[4]), .ZN(n1) );
  INVX0 U229 ( .INP(SH[3]), .ZN(n17) );
  INVX0 U230 ( .INP(SH[2]), .ZN(n58) );
  INVX0 U231 ( .INP(SH[1]), .ZN(n95) );
  AND2X1 U232 ( .IN1(n56), .IN2(n1), .Q(B[31]) );
  AND2X1 U233 ( .IN1(n55), .IN2(n1), .Q(B[30]) );
  AND2X1 U234 ( .IN1(A[32]), .IN2(n130), .Q(n163) );
  INVX0 U235 ( .INP(SH[0]), .ZN(n130) );
endmodule


module thumb_DW_rightsh_3 ( A, DATA_TC, SH, B );
  input [32:0] A;
  input [7:0] SH;
  output [32:0] B;
  input DATA_TC;
  wire   n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n44, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n81, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n118, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n155, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n191, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n307;

  AND2X1 U4 ( .IN1(n41), .IN2(n307), .Q(B[32]) );
  AND2X1 U5 ( .IN1(n40), .IN2(n307), .Q(B[31]) );
  AND2X1 U6 ( .IN1(n39), .IN2(n307), .Q(B[30]) );
  AND2X1 U7 ( .IN1(n38), .IN2(n307), .Q(B[29]) );
  AND2X1 U8 ( .IN1(n37), .IN2(n307), .Q(B[28]) );
  AND2X1 U9 ( .IN1(n36), .IN2(n307), .Q(B[27]) );
  AND2X1 U10 ( .IN1(n35), .IN2(n307), .Q(B[26]) );
  AND2X1 U11 ( .IN1(n34), .IN2(n307), .Q(B[25]) );
  AND2X1 U12 ( .IN1(n33), .IN2(n307), .Q(B[24]) );
  AND2X1 U13 ( .IN1(n32), .IN2(n307), .Q(B[23]) );
  AND2X1 U14 ( .IN1(n31), .IN2(n307), .Q(B[22]) );
  AND2X1 U15 ( .IN1(n30), .IN2(n307), .Q(B[21]) );
  AND2X1 U16 ( .IN1(n29), .IN2(n307), .Q(B[20]) );
  AND2X1 U17 ( .IN1(n28), .IN2(n307), .Q(B[19]) );
  AND2X1 U18 ( .IN1(n27), .IN2(n307), .Q(B[18]) );
  AND2X1 U19 ( .IN1(n26), .IN2(n307), .Q(B[17]) );
  AND2X1 U20 ( .IN1(n25), .IN2(n307), .Q(B[16]) );
  AND2X1 U21 ( .IN1(n24), .IN2(n307), .Q(B[15]) );
  AND2X1 U22 ( .IN1(n23), .IN2(n307), .Q(B[14]) );
  AND2X1 U23 ( .IN1(n22), .IN2(n307), .Q(B[13]) );
  AND2X1 U24 ( .IN1(n21), .IN2(n307), .Q(B[12]) );
  AND2X1 U25 ( .IN1(n20), .IN2(n307), .Q(B[11]) );
  AND2X1 U26 ( .IN1(n19), .IN2(n307), .Q(B[10]) );
  AND2X1 U27 ( .IN1(n18), .IN2(n307), .Q(B[9]) );
  AND2X1 U28 ( .IN1(n17), .IN2(n307), .Q(B[8]) );
  AND2X1 U29 ( .IN1(n16), .IN2(n307), .Q(B[7]) );
  AND2X1 U30 ( .IN1(n15), .IN2(n307), .Q(B[6]) );
  AND2X1 U31 ( .IN1(n14), .IN2(n307), .Q(B[5]) );
  AND2X1 U32 ( .IN1(n13), .IN2(n307), .Q(B[4]) );
  AND2X1 U33 ( .IN1(n12), .IN2(n307), .Q(B[3]) );
  AND2X1 U34 ( .IN1(n11), .IN2(n307), .Q(B[2]) );
  AND2X1 U35 ( .IN1(n10), .IN2(n307), .Q(B[1]) );
  AND2X1 U36 ( .IN1(n9), .IN2(n307), .Q(B[0]) );
  AND2X1 U41 ( .IN1(n78), .IN2(n7), .Q(n41) );
  AND2X1 U42 ( .IN1(n77), .IN2(n7), .Q(n40) );
  AND2X1 U43 ( .IN1(n76), .IN2(n7), .Q(n39) );
  AND2X1 U44 ( .IN1(n75), .IN2(n7), .Q(n38) );
  AND2X1 U45 ( .IN1(n74), .IN2(n7), .Q(n37) );
  AND2X1 U46 ( .IN1(n73), .IN2(n7), .Q(n36) );
  AND2X1 U47 ( .IN1(n72), .IN2(n7), .Q(n35) );
  AND2X1 U48 ( .IN1(n71), .IN2(n7), .Q(n34) );
  AND2X1 U49 ( .IN1(n70), .IN2(n7), .Q(n33) );
  AND2X1 U50 ( .IN1(n69), .IN2(n7), .Q(n32) );
  AND2X1 U51 ( .IN1(n68), .IN2(n7), .Q(n31) );
  AND2X1 U52 ( .IN1(n67), .IN2(n7), .Q(n30) );
  AND2X1 U53 ( .IN1(n66), .IN2(n7), .Q(n29) );
  AND2X1 U54 ( .IN1(n65), .IN2(n7), .Q(n28) );
  AND2X1 U55 ( .IN1(n64), .IN2(n7), .Q(n27) );
  AND2X1 U56 ( .IN1(n63), .IN2(n7), .Q(n26) );
  AND2X1 U57 ( .IN1(n62), .IN2(n7), .Q(n25) );
  AND2X1 U58 ( .IN1(n61), .IN2(n7), .Q(n24) );
  AND2X1 U59 ( .IN1(n60), .IN2(n7), .Q(n23) );
  AND2X1 U60 ( .IN1(n59), .IN2(n7), .Q(n22) );
  AND2X1 U61 ( .IN1(n58), .IN2(n7), .Q(n21) );
  AND2X1 U62 ( .IN1(n57), .IN2(n7), .Q(n20) );
  AND2X1 U63 ( .IN1(n56), .IN2(n7), .Q(n19) );
  AND2X1 U64 ( .IN1(n55), .IN2(n7), .Q(n18) );
  AND2X1 U65 ( .IN1(n54), .IN2(n7), .Q(n17) );
  AND2X1 U66 ( .IN1(n53), .IN2(n7), .Q(n16) );
  AND2X1 U67 ( .IN1(n52), .IN2(n7), .Q(n15) );
  AND2X1 U68 ( .IN1(n51), .IN2(n7), .Q(n14) );
  AND2X1 U69 ( .IN1(n50), .IN2(n7), .Q(n13) );
  AND2X1 U70 ( .IN1(n49), .IN2(n7), .Q(n12) );
  AND2X1 U71 ( .IN1(n48), .IN2(n7), .Q(n11) );
  AND2X1 U72 ( .IN1(n47), .IN2(n7), .Q(n10) );
  AO22X1 U73 ( .IN1(SH[5]), .IN2(n78), .IN3(n46), .IN4(n7), .Q(n9) );
  AND2X1 U78 ( .IN1(n115), .IN2(n44), .Q(n78) );
  AND2X1 U79 ( .IN1(n114), .IN2(n44), .Q(n77) );
  AND2X1 U80 ( .IN1(n113), .IN2(n44), .Q(n76) );
  AND2X1 U81 ( .IN1(n112), .IN2(n44), .Q(n75) );
  AND2X1 U82 ( .IN1(n111), .IN2(n44), .Q(n74) );
  AND2X1 U83 ( .IN1(n110), .IN2(n44), .Q(n73) );
  AND2X1 U84 ( .IN1(n109), .IN2(n44), .Q(n72) );
  AND2X1 U85 ( .IN1(n108), .IN2(n44), .Q(n71) );
  AND2X1 U86 ( .IN1(n107), .IN2(n44), .Q(n70) );
  AND2X1 U87 ( .IN1(n106), .IN2(n44), .Q(n69) );
  AND2X1 U88 ( .IN1(n105), .IN2(n44), .Q(n68) );
  AND2X1 U89 ( .IN1(n104), .IN2(n44), .Q(n67) );
  AND2X1 U90 ( .IN1(n103), .IN2(n44), .Q(n66) );
  AND2X1 U91 ( .IN1(n102), .IN2(n44), .Q(n65) );
  AND2X1 U92 ( .IN1(n101), .IN2(n44), .Q(n64) );
  AND2X1 U93 ( .IN1(n100), .IN2(n44), .Q(n63) );
  AO22X1 U94 ( .IN1(SH[4]), .IN2(n115), .IN3(n99), .IN4(n44), .Q(n62) );
  AO22X1 U95 ( .IN1(SH[4]), .IN2(n114), .IN3(n98), .IN4(n44), .Q(n61) );
  AO22X1 U96 ( .IN1(SH[4]), .IN2(n113), .IN3(n97), .IN4(n44), .Q(n60) );
  AO22X1 U97 ( .IN1(SH[4]), .IN2(n112), .IN3(n96), .IN4(n44), .Q(n59) );
  AO22X1 U98 ( .IN1(SH[4]), .IN2(n111), .IN3(n95), .IN4(n44), .Q(n58) );
  AO22X1 U99 ( .IN1(SH[4]), .IN2(n110), .IN3(n94), .IN4(n44), .Q(n57) );
  AO22X1 U100 ( .IN1(SH[4]), .IN2(n109), .IN3(n93), .IN4(n44), .Q(n56) );
  AO22X1 U101 ( .IN1(SH[4]), .IN2(n108), .IN3(n92), .IN4(n44), .Q(n55) );
  AO22X1 U102 ( .IN1(SH[4]), .IN2(n107), .IN3(n91), .IN4(n44), .Q(n54) );
  AO22X1 U103 ( .IN1(SH[4]), .IN2(n106), .IN3(n90), .IN4(n44), .Q(n53) );
  AO22X1 U104 ( .IN1(SH[4]), .IN2(n105), .IN3(n89), .IN4(n44), .Q(n52) );
  AO22X1 U105 ( .IN1(SH[4]), .IN2(n104), .IN3(n88), .IN4(n44), .Q(n51) );
  AO22X1 U106 ( .IN1(SH[4]), .IN2(n103), .IN3(n87), .IN4(n44), .Q(n50) );
  AO22X1 U107 ( .IN1(SH[4]), .IN2(n102), .IN3(n86), .IN4(n44), .Q(n49) );
  AO22X1 U108 ( .IN1(SH[4]), .IN2(n101), .IN3(n85), .IN4(n44), .Q(n48) );
  AO22X1 U109 ( .IN1(SH[4]), .IN2(n100), .IN3(n84), .IN4(n44), .Q(n47) );
  AO22X1 U110 ( .IN1(n44), .IN2(n83), .IN3(n99), .IN4(SH[4]), .Q(n46) );
  AND2X1 U115 ( .IN1(n152), .IN2(n81), .Q(n115) );
  AND2X1 U116 ( .IN1(n151), .IN2(n81), .Q(n114) );
  AND2X1 U117 ( .IN1(n150), .IN2(n81), .Q(n113) );
  AND2X1 U118 ( .IN1(n149), .IN2(n81), .Q(n112) );
  AND2X1 U119 ( .IN1(n148), .IN2(n81), .Q(n111) );
  AND2X1 U120 ( .IN1(n147), .IN2(n81), .Q(n110) );
  AND2X1 U121 ( .IN1(n146), .IN2(n81), .Q(n109) );
  AND2X1 U122 ( .IN1(n145), .IN2(n81), .Q(n108) );
  AO22X1 U123 ( .IN1(SH[3]), .IN2(n152), .IN3(n144), .IN4(n81), .Q(n107) );
  AO22X1 U124 ( .IN1(SH[3]), .IN2(n151), .IN3(n143), .IN4(n81), .Q(n106) );
  AO22X1 U125 ( .IN1(SH[3]), .IN2(n150), .IN3(n142), .IN4(n81), .Q(n105) );
  AO22X1 U126 ( .IN1(SH[3]), .IN2(n149), .IN3(n141), .IN4(n81), .Q(n104) );
  AO22X1 U127 ( .IN1(SH[3]), .IN2(n148), .IN3(n140), .IN4(n81), .Q(n103) );
  AO22X1 U128 ( .IN1(SH[3]), .IN2(n147), .IN3(n139), .IN4(n81), .Q(n102) );
  AO22X1 U129 ( .IN1(SH[3]), .IN2(n146), .IN3(n138), .IN4(n81), .Q(n101) );
  AO22X1 U130 ( .IN1(SH[3]), .IN2(n145), .IN3(n137), .IN4(n81), .Q(n100) );
  AO22X1 U131 ( .IN1(SH[3]), .IN2(n144), .IN3(n136), .IN4(n81), .Q(n99) );
  AO22X1 U132 ( .IN1(SH[3]), .IN2(n143), .IN3(n135), .IN4(n81), .Q(n98) );
  AO22X1 U133 ( .IN1(SH[3]), .IN2(n142), .IN3(n134), .IN4(n81), .Q(n97) );
  AO22X1 U134 ( .IN1(SH[3]), .IN2(n141), .IN3(n133), .IN4(n81), .Q(n96) );
  AO22X1 U135 ( .IN1(SH[3]), .IN2(n140), .IN3(n132), .IN4(n81), .Q(n95) );
  AO22X1 U136 ( .IN1(SH[3]), .IN2(n139), .IN3(n131), .IN4(n81), .Q(n94) );
  AO22X1 U137 ( .IN1(SH[3]), .IN2(n138), .IN3(n130), .IN4(n81), .Q(n93) );
  AO22X1 U138 ( .IN1(SH[3]), .IN2(n137), .IN3(n129), .IN4(n81), .Q(n92) );
  AO22X1 U139 ( .IN1(SH[3]), .IN2(n136), .IN3(n128), .IN4(n81), .Q(n91) );
  AO22X1 U140 ( .IN1(SH[3]), .IN2(n135), .IN3(n127), .IN4(n81), .Q(n90) );
  AO22X1 U141 ( .IN1(SH[3]), .IN2(n134), .IN3(n126), .IN4(n81), .Q(n89) );
  AO22X1 U142 ( .IN1(SH[3]), .IN2(n133), .IN3(n125), .IN4(n81), .Q(n88) );
  AO22X1 U143 ( .IN1(SH[3]), .IN2(n132), .IN3(n124), .IN4(n81), .Q(n87) );
  AO22X1 U144 ( .IN1(SH[3]), .IN2(n131), .IN3(n123), .IN4(n81), .Q(n86) );
  AO22X1 U145 ( .IN1(SH[3]), .IN2(n130), .IN3(n122), .IN4(n81), .Q(n85) );
  AO22X1 U146 ( .IN1(SH[3]), .IN2(n129), .IN3(n121), .IN4(n81), .Q(n84) );
  AO22X1 U147 ( .IN1(n81), .IN2(n120), .IN3(n128), .IN4(SH[3]), .Q(n83) );
  AND2X1 U152 ( .IN1(n189), .IN2(n118), .Q(n152) );
  AND2X1 U153 ( .IN1(n188), .IN2(n118), .Q(n151) );
  AND2X1 U154 ( .IN1(n187), .IN2(n118), .Q(n150) );
  AND2X1 U155 ( .IN1(n186), .IN2(n118), .Q(n149) );
  AO22X1 U156 ( .IN1(SH[2]), .IN2(n189), .IN3(n185), .IN4(n118), .Q(n148) );
  AO22X1 U157 ( .IN1(SH[2]), .IN2(n188), .IN3(n184), .IN4(n118), .Q(n147) );
  AO22X1 U158 ( .IN1(SH[2]), .IN2(n187), .IN3(n183), .IN4(n118), .Q(n146) );
  AO22X1 U159 ( .IN1(SH[2]), .IN2(n186), .IN3(n182), .IN4(n118), .Q(n145) );
  AO22X1 U160 ( .IN1(SH[2]), .IN2(n185), .IN3(n181), .IN4(n118), .Q(n144) );
  AO22X1 U161 ( .IN1(SH[2]), .IN2(n184), .IN3(n180), .IN4(n118), .Q(n143) );
  AO22X1 U162 ( .IN1(SH[2]), .IN2(n183), .IN3(n179), .IN4(n118), .Q(n142) );
  AO22X1 U163 ( .IN1(SH[2]), .IN2(n182), .IN3(n178), .IN4(n118), .Q(n141) );
  AO22X1 U164 ( .IN1(SH[2]), .IN2(n181), .IN3(n177), .IN4(n118), .Q(n140) );
  AO22X1 U165 ( .IN1(SH[2]), .IN2(n180), .IN3(n176), .IN4(n118), .Q(n139) );
  AO22X1 U166 ( .IN1(SH[2]), .IN2(n179), .IN3(n175), .IN4(n118), .Q(n138) );
  AO22X1 U167 ( .IN1(SH[2]), .IN2(n178), .IN3(n174), .IN4(n118), .Q(n137) );
  AO22X1 U168 ( .IN1(SH[2]), .IN2(n177), .IN3(n173), .IN4(n118), .Q(n136) );
  AO22X1 U169 ( .IN1(SH[2]), .IN2(n176), .IN3(n172), .IN4(n118), .Q(n135) );
  AO22X1 U170 ( .IN1(SH[2]), .IN2(n175), .IN3(n171), .IN4(n118), .Q(n134) );
  AO22X1 U171 ( .IN1(SH[2]), .IN2(n174), .IN3(n170), .IN4(n118), .Q(n133) );
  AO22X1 U172 ( .IN1(SH[2]), .IN2(n173), .IN3(n169), .IN4(n118), .Q(n132) );
  AO22X1 U173 ( .IN1(SH[2]), .IN2(n172), .IN3(n168), .IN4(n118), .Q(n131) );
  AO22X1 U174 ( .IN1(SH[2]), .IN2(n171), .IN3(n167), .IN4(n118), .Q(n130) );
  AO22X1 U175 ( .IN1(SH[2]), .IN2(n170), .IN3(n166), .IN4(n118), .Q(n129) );
  AO22X1 U176 ( .IN1(SH[2]), .IN2(n169), .IN3(n165), .IN4(n118), .Q(n128) );
  AO22X1 U177 ( .IN1(SH[2]), .IN2(n168), .IN3(n164), .IN4(n118), .Q(n127) );
  AO22X1 U178 ( .IN1(SH[2]), .IN2(n167), .IN3(n163), .IN4(n118), .Q(n126) );
  AO22X1 U179 ( .IN1(SH[2]), .IN2(n166), .IN3(n162), .IN4(n118), .Q(n125) );
  AO22X1 U180 ( .IN1(SH[2]), .IN2(n165), .IN3(n161), .IN4(n118), .Q(n124) );
  AO22X1 U181 ( .IN1(SH[2]), .IN2(n164), .IN3(n160), .IN4(n118), .Q(n123) );
  AO22X1 U182 ( .IN1(SH[2]), .IN2(n163), .IN3(n159), .IN4(n118), .Q(n122) );
  AO22X1 U183 ( .IN1(SH[2]), .IN2(n162), .IN3(n158), .IN4(n118), .Q(n121) );
  AO22X1 U184 ( .IN1(n118), .IN2(n157), .IN3(n161), .IN4(SH[2]), .Q(n120) );
  AND2X1 U189 ( .IN1(n225), .IN2(n155), .Q(n189) );
  AND2X1 U190 ( .IN1(n224), .IN2(n155), .Q(n188) );
  AO22X1 U191 ( .IN1(SH[1]), .IN2(n225), .IN3(n223), .IN4(n155), .Q(n187) );
  AO22X1 U192 ( .IN1(SH[1]), .IN2(n224), .IN3(n222), .IN4(n155), .Q(n186) );
  AO22X1 U193 ( .IN1(SH[1]), .IN2(n223), .IN3(n221), .IN4(n155), .Q(n185) );
  AO22X1 U194 ( .IN1(SH[1]), .IN2(n222), .IN3(n220), .IN4(n155), .Q(n184) );
  AO22X1 U195 ( .IN1(SH[1]), .IN2(n221), .IN3(n219), .IN4(n155), .Q(n183) );
  AO22X1 U196 ( .IN1(SH[1]), .IN2(n220), .IN3(n218), .IN4(n155), .Q(n182) );
  AO22X1 U197 ( .IN1(SH[1]), .IN2(n219), .IN3(n217), .IN4(n155), .Q(n181) );
  AO22X1 U198 ( .IN1(SH[1]), .IN2(n218), .IN3(n216), .IN4(n155), .Q(n180) );
  AO22X1 U199 ( .IN1(SH[1]), .IN2(n217), .IN3(n215), .IN4(n155), .Q(n179) );
  AO22X1 U200 ( .IN1(SH[1]), .IN2(n216), .IN3(n214), .IN4(n155), .Q(n178) );
  AO22X1 U201 ( .IN1(SH[1]), .IN2(n215), .IN3(n213), .IN4(n155), .Q(n177) );
  AO22X1 U202 ( .IN1(SH[1]), .IN2(n214), .IN3(n212), .IN4(n155), .Q(n176) );
  AO22X1 U203 ( .IN1(SH[1]), .IN2(n213), .IN3(n211), .IN4(n155), .Q(n175) );
  AO22X1 U204 ( .IN1(SH[1]), .IN2(n212), .IN3(n210), .IN4(n155), .Q(n174) );
  AO22X1 U205 ( .IN1(SH[1]), .IN2(n211), .IN3(n209), .IN4(n155), .Q(n173) );
  AO22X1 U206 ( .IN1(SH[1]), .IN2(n210), .IN3(n208), .IN4(n155), .Q(n172) );
  AO22X1 U207 ( .IN1(SH[1]), .IN2(n209), .IN3(n207), .IN4(n155), .Q(n171) );
  AO22X1 U208 ( .IN1(SH[1]), .IN2(n208), .IN3(n206), .IN4(n155), .Q(n170) );
  AO22X1 U209 ( .IN1(SH[1]), .IN2(n207), .IN3(n205), .IN4(n155), .Q(n169) );
  AO22X1 U210 ( .IN1(SH[1]), .IN2(n206), .IN3(n204), .IN4(n155), .Q(n168) );
  AO22X1 U211 ( .IN1(SH[1]), .IN2(n205), .IN3(n203), .IN4(n155), .Q(n167) );
  AO22X1 U212 ( .IN1(SH[1]), .IN2(n204), .IN3(n202), .IN4(n155), .Q(n166) );
  AO22X1 U213 ( .IN1(SH[1]), .IN2(n203), .IN3(n201), .IN4(n155), .Q(n165) );
  AO22X1 U214 ( .IN1(SH[1]), .IN2(n202), .IN3(n200), .IN4(n155), .Q(n164) );
  AO22X1 U215 ( .IN1(SH[1]), .IN2(n201), .IN3(n199), .IN4(n155), .Q(n163) );
  AO22X1 U216 ( .IN1(SH[1]), .IN2(n200), .IN3(n198), .IN4(n155), .Q(n162) );
  AO22X1 U217 ( .IN1(SH[1]), .IN2(n199), .IN3(n197), .IN4(n155), .Q(n161) );
  AO22X1 U218 ( .IN1(SH[1]), .IN2(n198), .IN3(n196), .IN4(n155), .Q(n160) );
  AO22X1 U219 ( .IN1(SH[1]), .IN2(n197), .IN3(n195), .IN4(n155), .Q(n159) );
  AO22X1 U220 ( .IN1(SH[1]), .IN2(n196), .IN3(n194), .IN4(n155), .Q(n158) );
  AO22X1 U221 ( .IN1(n193), .IN2(n155), .IN3(n195), .IN4(SH[1]), .Q(n157) );
  AND2X1 U225 ( .IN1(n191), .IN2(A[32]), .Q(n225) );
  AO22X1 U226 ( .IN1(A[32]), .IN2(SH[0]), .IN3(n191), .IN4(A[31]), .Q(n224) );
  AO22X1 U227 ( .IN1(A[31]), .IN2(SH[0]), .IN3(n191), .IN4(A[30]), .Q(n223) );
  AO22X1 U228 ( .IN1(A[30]), .IN2(SH[0]), .IN3(n191), .IN4(A[29]), .Q(n222) );
  AO22X1 U229 ( .IN1(A[29]), .IN2(SH[0]), .IN3(n191), .IN4(A[28]), .Q(n221) );
  AO22X1 U230 ( .IN1(A[28]), .IN2(SH[0]), .IN3(n191), .IN4(A[27]), .Q(n220) );
  AO22X1 U231 ( .IN1(A[27]), .IN2(SH[0]), .IN3(n191), .IN4(A[26]), .Q(n219) );
  AO22X1 U232 ( .IN1(A[26]), .IN2(SH[0]), .IN3(n191), .IN4(A[25]), .Q(n218) );
  AO22X1 U233 ( .IN1(A[25]), .IN2(SH[0]), .IN3(n191), .IN4(A[24]), .Q(n217) );
  AO22X1 U234 ( .IN1(A[24]), .IN2(SH[0]), .IN3(n191), .IN4(A[23]), .Q(n216) );
  AO22X1 U235 ( .IN1(A[23]), .IN2(SH[0]), .IN3(n191), .IN4(A[22]), .Q(n215) );
  AO22X1 U236 ( .IN1(A[22]), .IN2(SH[0]), .IN3(n191), .IN4(A[21]), .Q(n214) );
  AO22X1 U237 ( .IN1(A[21]), .IN2(SH[0]), .IN3(n191), .IN4(A[20]), .Q(n213) );
  AO22X1 U238 ( .IN1(A[20]), .IN2(SH[0]), .IN3(n191), .IN4(A[19]), .Q(n212) );
  AO22X1 U239 ( .IN1(A[19]), .IN2(SH[0]), .IN3(n191), .IN4(A[18]), .Q(n211) );
  AO22X1 U240 ( .IN1(A[18]), .IN2(SH[0]), .IN3(n191), .IN4(A[17]), .Q(n210) );
  AO22X1 U241 ( .IN1(A[17]), .IN2(SH[0]), .IN3(n191), .IN4(A[16]), .Q(n209) );
  AO22X1 U242 ( .IN1(A[16]), .IN2(SH[0]), .IN3(n191), .IN4(A[15]), .Q(n208) );
  AO22X1 U243 ( .IN1(A[15]), .IN2(SH[0]), .IN3(n191), .IN4(A[14]), .Q(n207) );
  AO22X1 U244 ( .IN1(A[14]), .IN2(SH[0]), .IN3(n191), .IN4(A[13]), .Q(n206) );
  AO22X1 U245 ( .IN1(A[13]), .IN2(SH[0]), .IN3(n191), .IN4(A[12]), .Q(n205) );
  AO22X1 U246 ( .IN1(A[12]), .IN2(SH[0]), .IN3(n191), .IN4(A[11]), .Q(n204) );
  AO22X1 U247 ( .IN1(A[11]), .IN2(SH[0]), .IN3(n191), .IN4(A[10]), .Q(n203) );
  AO22X1 U248 ( .IN1(A[10]), .IN2(SH[0]), .IN3(n191), .IN4(A[9]), .Q(n202) );
  AO22X1 U249 ( .IN1(A[9]), .IN2(SH[0]), .IN3(n191), .IN4(A[8]), .Q(n201) );
  AO22X1 U250 ( .IN1(A[8]), .IN2(SH[0]), .IN3(n191), .IN4(A[7]), .Q(n200) );
  AO22X1 U251 ( .IN1(A[7]), .IN2(SH[0]), .IN3(n191), .IN4(A[6]), .Q(n199) );
  AO22X1 U252 ( .IN1(A[6]), .IN2(SH[0]), .IN3(n191), .IN4(A[5]), .Q(n198) );
  AO22X1 U253 ( .IN1(A[5]), .IN2(SH[0]), .IN3(n191), .IN4(A[4]), .Q(n197) );
  AO22X1 U254 ( .IN1(A[4]), .IN2(SH[0]), .IN3(n191), .IN4(A[3]), .Q(n196) );
  AO22X1 U255 ( .IN1(A[3]), .IN2(SH[0]), .IN3(n191), .IN4(A[2]), .Q(n195) );
  AO22X1 U256 ( .IN1(A[2]), .IN2(SH[0]), .IN3(n191), .IN4(A[1]), .Q(n194) );
  AND2X1 U257 ( .IN1(SH[0]), .IN2(A[1]), .Q(n193) );
  INVX0 U263 ( .INP(SH[1]), .ZN(n155) );
  INVX0 U264 ( .INP(SH[2]), .ZN(n118) );
  INVX0 U265 ( .INP(SH[0]), .ZN(n191) );
  INVX0 U266 ( .INP(SH[3]), .ZN(n81) );
  INVX0 U267 ( .INP(SH[4]), .ZN(n44) );
  INVX0 U268 ( .INP(SH[5]), .ZN(n7) );
  NOR2X0 U269 ( .IN1(SH[7]), .IN2(SH[6]), .QN(n307) );
endmodule


module thumb_DW_leftsh_3 ( A, SH, B );
  input [32:0] A;
  input [7:0] SH;
  output [32:0] B;
  wire   n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n44, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n81, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n118, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n155, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n191, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n306;

  AND2X1 U4 ( .IN1(n41), .IN2(n306), .Q(B[32]) );
  AND2X1 U5 ( .IN1(n40), .IN2(n306), .Q(B[31]) );
  AND2X1 U6 ( .IN1(n39), .IN2(n306), .Q(B[30]) );
  AND2X1 U7 ( .IN1(n38), .IN2(n306), .Q(B[29]) );
  AND2X1 U8 ( .IN1(n37), .IN2(n306), .Q(B[28]) );
  AND2X1 U9 ( .IN1(n36), .IN2(n306), .Q(B[27]) );
  AND2X1 U10 ( .IN1(n35), .IN2(n306), .Q(B[26]) );
  AND2X1 U11 ( .IN1(n34), .IN2(n306), .Q(B[25]) );
  AND2X1 U12 ( .IN1(n33), .IN2(n306), .Q(B[24]) );
  AND2X1 U13 ( .IN1(n32), .IN2(n306), .Q(B[23]) );
  AND2X1 U14 ( .IN1(n31), .IN2(n306), .Q(B[22]) );
  AND2X1 U15 ( .IN1(n30), .IN2(n306), .Q(B[21]) );
  AND2X1 U16 ( .IN1(n29), .IN2(n306), .Q(B[20]) );
  AND2X1 U17 ( .IN1(n28), .IN2(n306), .Q(B[19]) );
  AND2X1 U18 ( .IN1(n27), .IN2(n306), .Q(B[18]) );
  AND2X1 U19 ( .IN1(n26), .IN2(n306), .Q(B[17]) );
  AND2X1 U20 ( .IN1(n25), .IN2(n306), .Q(B[16]) );
  AND2X1 U21 ( .IN1(n24), .IN2(n306), .Q(B[15]) );
  AND2X1 U22 ( .IN1(n23), .IN2(n306), .Q(B[14]) );
  AND2X1 U23 ( .IN1(n22), .IN2(n306), .Q(B[13]) );
  AND2X1 U24 ( .IN1(n21), .IN2(n306), .Q(B[12]) );
  AND2X1 U25 ( .IN1(n20), .IN2(n306), .Q(B[11]) );
  AND2X1 U26 ( .IN1(n19), .IN2(n306), .Q(B[10]) );
  AND2X1 U27 ( .IN1(n18), .IN2(n306), .Q(B[9]) );
  AND2X1 U28 ( .IN1(n17), .IN2(n306), .Q(B[8]) );
  AND2X1 U29 ( .IN1(n16), .IN2(n306), .Q(B[7]) );
  AND2X1 U30 ( .IN1(n15), .IN2(n306), .Q(B[6]) );
  AND2X1 U31 ( .IN1(n14), .IN2(n306), .Q(B[5]) );
  AND2X1 U32 ( .IN1(n13), .IN2(n306), .Q(B[4]) );
  AND2X1 U33 ( .IN1(n12), .IN2(n306), .Q(B[3]) );
  AND2X1 U34 ( .IN1(n11), .IN2(n306), .Q(B[2]) );
  AND2X1 U35 ( .IN1(n10), .IN2(n306), .Q(B[1]) );
  AND2X1 U36 ( .IN1(n9), .IN2(n306), .Q(B[0]) );
  AO22X1 U41 ( .IN1(SH[5]), .IN2(n46), .IN3(n78), .IN4(n7), .Q(n41) );
  AND2X1 U42 ( .IN1(n77), .IN2(n7), .Q(n40) );
  AND2X1 U43 ( .IN1(n76), .IN2(n7), .Q(n39) );
  AND2X1 U44 ( .IN1(n75), .IN2(n7), .Q(n38) );
  AND2X1 U45 ( .IN1(n74), .IN2(n7), .Q(n37) );
  AND2X1 U46 ( .IN1(n73), .IN2(n7), .Q(n36) );
  AND2X1 U47 ( .IN1(n72), .IN2(n7), .Q(n35) );
  AND2X1 U48 ( .IN1(n71), .IN2(n7), .Q(n34) );
  AND2X1 U49 ( .IN1(n70), .IN2(n7), .Q(n33) );
  AND2X1 U50 ( .IN1(n69), .IN2(n7), .Q(n32) );
  AND2X1 U51 ( .IN1(n68), .IN2(n7), .Q(n31) );
  AND2X1 U52 ( .IN1(n67), .IN2(n7), .Q(n30) );
  AND2X1 U53 ( .IN1(n66), .IN2(n7), .Q(n29) );
  AND2X1 U54 ( .IN1(n65), .IN2(n7), .Q(n28) );
  AND2X1 U55 ( .IN1(n64), .IN2(n7), .Q(n27) );
  AND2X1 U56 ( .IN1(n63), .IN2(n7), .Q(n26) );
  AND2X1 U57 ( .IN1(n62), .IN2(n7), .Q(n25) );
  AND2X1 U58 ( .IN1(n61), .IN2(n7), .Q(n24) );
  AND2X1 U59 ( .IN1(n60), .IN2(n7), .Q(n23) );
  AND2X1 U60 ( .IN1(n59), .IN2(n7), .Q(n22) );
  AND2X1 U61 ( .IN1(n58), .IN2(n7), .Q(n21) );
  AND2X1 U62 ( .IN1(n57), .IN2(n7), .Q(n20) );
  AND2X1 U63 ( .IN1(n56), .IN2(n7), .Q(n19) );
  AND2X1 U64 ( .IN1(n55), .IN2(n7), .Q(n18) );
  AND2X1 U65 ( .IN1(n54), .IN2(n7), .Q(n17) );
  AND2X1 U66 ( .IN1(n53), .IN2(n7), .Q(n16) );
  AND2X1 U67 ( .IN1(n52), .IN2(n7), .Q(n15) );
  AND2X1 U68 ( .IN1(n51), .IN2(n7), .Q(n14) );
  AND2X1 U69 ( .IN1(n50), .IN2(n7), .Q(n13) );
  AND2X1 U70 ( .IN1(n49), .IN2(n7), .Q(n12) );
  AND2X1 U71 ( .IN1(n48), .IN2(n7), .Q(n11) );
  AND2X1 U72 ( .IN1(n47), .IN2(n7), .Q(n10) );
  AND2X1 U73 ( .IN1(n46), .IN2(n7), .Q(n9) );
  AO22X1 U78 ( .IN1(n44), .IN2(n115), .IN3(n99), .IN4(SH[4]), .Q(n78) );
  AO22X1 U79 ( .IN1(SH[4]), .IN2(n98), .IN3(n114), .IN4(n44), .Q(n77) );
  AO22X1 U80 ( .IN1(SH[4]), .IN2(n97), .IN3(n113), .IN4(n44), .Q(n76) );
  AO22X1 U81 ( .IN1(SH[4]), .IN2(n96), .IN3(n112), .IN4(n44), .Q(n75) );
  AO22X1 U82 ( .IN1(SH[4]), .IN2(n95), .IN3(n111), .IN4(n44), .Q(n74) );
  AO22X1 U83 ( .IN1(SH[4]), .IN2(n94), .IN3(n110), .IN4(n44), .Q(n73) );
  AO22X1 U84 ( .IN1(SH[4]), .IN2(n93), .IN3(n109), .IN4(n44), .Q(n72) );
  AO22X1 U85 ( .IN1(SH[4]), .IN2(n92), .IN3(n108), .IN4(n44), .Q(n71) );
  AO22X1 U86 ( .IN1(SH[4]), .IN2(n91), .IN3(n107), .IN4(n44), .Q(n70) );
  AO22X1 U87 ( .IN1(SH[4]), .IN2(n90), .IN3(n106), .IN4(n44), .Q(n69) );
  AO22X1 U88 ( .IN1(SH[4]), .IN2(n89), .IN3(n105), .IN4(n44), .Q(n68) );
  AO22X1 U89 ( .IN1(SH[4]), .IN2(n88), .IN3(n104), .IN4(n44), .Q(n67) );
  AO22X1 U90 ( .IN1(SH[4]), .IN2(n87), .IN3(n103), .IN4(n44), .Q(n66) );
  AO22X1 U91 ( .IN1(SH[4]), .IN2(n86), .IN3(n102), .IN4(n44), .Q(n65) );
  AO22X1 U92 ( .IN1(SH[4]), .IN2(n85), .IN3(n101), .IN4(n44), .Q(n64) );
  AO22X1 U93 ( .IN1(SH[4]), .IN2(n84), .IN3(n100), .IN4(n44), .Q(n63) );
  AO22X1 U94 ( .IN1(SH[4]), .IN2(n83), .IN3(n99), .IN4(n44), .Q(n62) );
  AND2X1 U95 ( .IN1(n98), .IN2(n44), .Q(n61) );
  AND2X1 U96 ( .IN1(n97), .IN2(n44), .Q(n60) );
  AND2X1 U97 ( .IN1(n96), .IN2(n44), .Q(n59) );
  AND2X1 U98 ( .IN1(n95), .IN2(n44), .Q(n58) );
  AND2X1 U99 ( .IN1(n94), .IN2(n44), .Q(n57) );
  AND2X1 U100 ( .IN1(n93), .IN2(n44), .Q(n56) );
  AND2X1 U101 ( .IN1(n92), .IN2(n44), .Q(n55) );
  AND2X1 U102 ( .IN1(n91), .IN2(n44), .Q(n54) );
  AND2X1 U103 ( .IN1(n90), .IN2(n44), .Q(n53) );
  AND2X1 U104 ( .IN1(n89), .IN2(n44), .Q(n52) );
  AND2X1 U105 ( .IN1(n88), .IN2(n44), .Q(n51) );
  AND2X1 U106 ( .IN1(n87), .IN2(n44), .Q(n50) );
  AND2X1 U107 ( .IN1(n86), .IN2(n44), .Q(n49) );
  AND2X1 U108 ( .IN1(n85), .IN2(n44), .Q(n48) );
  AND2X1 U109 ( .IN1(n84), .IN2(n44), .Q(n47) );
  AND2X1 U110 ( .IN1(n83), .IN2(n44), .Q(n46) );
  AO22X1 U115 ( .IN1(n81), .IN2(n152), .IN3(n144), .IN4(SH[3]), .Q(n115) );
  AO22X1 U116 ( .IN1(SH[3]), .IN2(n143), .IN3(n151), .IN4(n81), .Q(n114) );
  AO22X1 U117 ( .IN1(SH[3]), .IN2(n142), .IN3(n150), .IN4(n81), .Q(n113) );
  AO22X1 U118 ( .IN1(SH[3]), .IN2(n141), .IN3(n149), .IN4(n81), .Q(n112) );
  AO22X1 U119 ( .IN1(SH[3]), .IN2(n140), .IN3(n148), .IN4(n81), .Q(n111) );
  AO22X1 U120 ( .IN1(SH[3]), .IN2(n139), .IN3(n147), .IN4(n81), .Q(n110) );
  AO22X1 U121 ( .IN1(SH[3]), .IN2(n138), .IN3(n146), .IN4(n81), .Q(n109) );
  AO22X1 U122 ( .IN1(SH[3]), .IN2(n137), .IN3(n145), .IN4(n81), .Q(n108) );
  AO22X1 U123 ( .IN1(SH[3]), .IN2(n136), .IN3(n144), .IN4(n81), .Q(n107) );
  AO22X1 U124 ( .IN1(SH[3]), .IN2(n135), .IN3(n143), .IN4(n81), .Q(n106) );
  AO22X1 U125 ( .IN1(SH[3]), .IN2(n134), .IN3(n142), .IN4(n81), .Q(n105) );
  AO22X1 U126 ( .IN1(SH[3]), .IN2(n133), .IN3(n141), .IN4(n81), .Q(n104) );
  AO22X1 U127 ( .IN1(SH[3]), .IN2(n132), .IN3(n140), .IN4(n81), .Q(n103) );
  AO22X1 U128 ( .IN1(SH[3]), .IN2(n131), .IN3(n139), .IN4(n81), .Q(n102) );
  AO22X1 U129 ( .IN1(SH[3]), .IN2(n130), .IN3(n138), .IN4(n81), .Q(n101) );
  AO22X1 U130 ( .IN1(SH[3]), .IN2(n129), .IN3(n137), .IN4(n81), .Q(n100) );
  AO22X1 U131 ( .IN1(SH[3]), .IN2(n128), .IN3(n136), .IN4(n81), .Q(n99) );
  AO22X1 U132 ( .IN1(SH[3]), .IN2(n127), .IN3(n135), .IN4(n81), .Q(n98) );
  AO22X1 U133 ( .IN1(SH[3]), .IN2(n126), .IN3(n134), .IN4(n81), .Q(n97) );
  AO22X1 U134 ( .IN1(SH[3]), .IN2(n125), .IN3(n133), .IN4(n81), .Q(n96) );
  AO22X1 U135 ( .IN1(SH[3]), .IN2(n124), .IN3(n132), .IN4(n81), .Q(n95) );
  AO22X1 U136 ( .IN1(SH[3]), .IN2(n123), .IN3(n131), .IN4(n81), .Q(n94) );
  AO22X1 U137 ( .IN1(SH[3]), .IN2(n122), .IN3(n130), .IN4(n81), .Q(n93) );
  AO22X1 U138 ( .IN1(SH[3]), .IN2(n121), .IN3(n129), .IN4(n81), .Q(n92) );
  AO22X1 U139 ( .IN1(SH[3]), .IN2(n120), .IN3(n128), .IN4(n81), .Q(n91) );
  AND2X1 U140 ( .IN1(n127), .IN2(n81), .Q(n90) );
  AND2X1 U141 ( .IN1(n126), .IN2(n81), .Q(n89) );
  AND2X1 U142 ( .IN1(n125), .IN2(n81), .Q(n88) );
  AND2X1 U143 ( .IN1(n124), .IN2(n81), .Q(n87) );
  AND2X1 U144 ( .IN1(n123), .IN2(n81), .Q(n86) );
  AND2X1 U145 ( .IN1(n122), .IN2(n81), .Q(n85) );
  AND2X1 U146 ( .IN1(n121), .IN2(n81), .Q(n84) );
  AND2X1 U147 ( .IN1(n120), .IN2(n81), .Q(n83) );
  AO22X1 U152 ( .IN1(n118), .IN2(n189), .IN3(n185), .IN4(SH[2]), .Q(n152) );
  AO22X1 U153 ( .IN1(SH[2]), .IN2(n184), .IN3(n188), .IN4(n118), .Q(n151) );
  AO22X1 U154 ( .IN1(SH[2]), .IN2(n183), .IN3(n187), .IN4(n118), .Q(n150) );
  AO22X1 U155 ( .IN1(SH[2]), .IN2(n182), .IN3(n186), .IN4(n118), .Q(n149) );
  AO22X1 U156 ( .IN1(SH[2]), .IN2(n181), .IN3(n185), .IN4(n118), .Q(n148) );
  AO22X1 U157 ( .IN1(SH[2]), .IN2(n180), .IN3(n184), .IN4(n118), .Q(n147) );
  AO22X1 U158 ( .IN1(SH[2]), .IN2(n179), .IN3(n183), .IN4(n118), .Q(n146) );
  AO22X1 U159 ( .IN1(SH[2]), .IN2(n178), .IN3(n182), .IN4(n118), .Q(n145) );
  AO22X1 U160 ( .IN1(SH[2]), .IN2(n177), .IN3(n181), .IN4(n118), .Q(n144) );
  AO22X1 U161 ( .IN1(SH[2]), .IN2(n176), .IN3(n180), .IN4(n118), .Q(n143) );
  AO22X1 U162 ( .IN1(SH[2]), .IN2(n175), .IN3(n179), .IN4(n118), .Q(n142) );
  AO22X1 U163 ( .IN1(SH[2]), .IN2(n174), .IN3(n178), .IN4(n118), .Q(n141) );
  AO22X1 U164 ( .IN1(SH[2]), .IN2(n173), .IN3(n177), .IN4(n118), .Q(n140) );
  AO22X1 U165 ( .IN1(SH[2]), .IN2(n172), .IN3(n176), .IN4(n118), .Q(n139) );
  AO22X1 U166 ( .IN1(SH[2]), .IN2(n171), .IN3(n175), .IN4(n118), .Q(n138) );
  AO22X1 U167 ( .IN1(SH[2]), .IN2(n170), .IN3(n174), .IN4(n118), .Q(n137) );
  AO22X1 U168 ( .IN1(SH[2]), .IN2(n169), .IN3(n173), .IN4(n118), .Q(n136) );
  AO22X1 U169 ( .IN1(SH[2]), .IN2(n168), .IN3(n172), .IN4(n118), .Q(n135) );
  AO22X1 U170 ( .IN1(SH[2]), .IN2(n167), .IN3(n171), .IN4(n118), .Q(n134) );
  AO22X1 U171 ( .IN1(SH[2]), .IN2(n166), .IN3(n170), .IN4(n118), .Q(n133) );
  AO22X1 U172 ( .IN1(SH[2]), .IN2(n165), .IN3(n169), .IN4(n118), .Q(n132) );
  AO22X1 U173 ( .IN1(SH[2]), .IN2(n164), .IN3(n168), .IN4(n118), .Q(n131) );
  AO22X1 U174 ( .IN1(SH[2]), .IN2(n163), .IN3(n167), .IN4(n118), .Q(n130) );
  AO22X1 U175 ( .IN1(SH[2]), .IN2(n162), .IN3(n166), .IN4(n118), .Q(n129) );
  AO22X1 U176 ( .IN1(SH[2]), .IN2(n161), .IN3(n165), .IN4(n118), .Q(n128) );
  AO22X1 U177 ( .IN1(SH[2]), .IN2(n160), .IN3(n164), .IN4(n118), .Q(n127) );
  AO22X1 U178 ( .IN1(SH[2]), .IN2(n159), .IN3(n163), .IN4(n118), .Q(n126) );
  AO22X1 U179 ( .IN1(SH[2]), .IN2(n158), .IN3(n162), .IN4(n118), .Q(n125) );
  AO22X1 U180 ( .IN1(SH[2]), .IN2(n157), .IN3(n161), .IN4(n118), .Q(n124) );
  AND2X1 U181 ( .IN1(n160), .IN2(n118), .Q(n123) );
  AND2X1 U182 ( .IN1(n159), .IN2(n118), .Q(n122) );
  AND2X1 U183 ( .IN1(n158), .IN2(n118), .Q(n121) );
  AND2X1 U184 ( .IN1(n157), .IN2(n118), .Q(n120) );
  AO22X1 U189 ( .IN1(n225), .IN2(n155), .IN3(n223), .IN4(SH[1]), .Q(n189) );
  AO22X1 U190 ( .IN1(SH[1]), .IN2(n222), .IN3(n224), .IN4(n155), .Q(n188) );
  AO22X1 U191 ( .IN1(SH[1]), .IN2(n221), .IN3(n223), .IN4(n155), .Q(n187) );
  AO22X1 U192 ( .IN1(SH[1]), .IN2(n220), .IN3(n222), .IN4(n155), .Q(n186) );
  AO22X1 U193 ( .IN1(SH[1]), .IN2(n219), .IN3(n221), .IN4(n155), .Q(n185) );
  AO22X1 U194 ( .IN1(SH[1]), .IN2(n218), .IN3(n220), .IN4(n155), .Q(n184) );
  AO22X1 U195 ( .IN1(SH[1]), .IN2(n217), .IN3(n219), .IN4(n155), .Q(n183) );
  AO22X1 U196 ( .IN1(SH[1]), .IN2(n216), .IN3(n218), .IN4(n155), .Q(n182) );
  AO22X1 U197 ( .IN1(SH[1]), .IN2(n215), .IN3(n217), .IN4(n155), .Q(n181) );
  AO22X1 U198 ( .IN1(SH[1]), .IN2(n214), .IN3(n216), .IN4(n155), .Q(n180) );
  AO22X1 U199 ( .IN1(SH[1]), .IN2(n213), .IN3(n215), .IN4(n155), .Q(n179) );
  AO22X1 U200 ( .IN1(SH[1]), .IN2(n212), .IN3(n214), .IN4(n155), .Q(n178) );
  AO22X1 U201 ( .IN1(SH[1]), .IN2(n211), .IN3(n213), .IN4(n155), .Q(n177) );
  AO22X1 U202 ( .IN1(SH[1]), .IN2(n210), .IN3(n212), .IN4(n155), .Q(n176) );
  AO22X1 U203 ( .IN1(SH[1]), .IN2(n209), .IN3(n211), .IN4(n155), .Q(n175) );
  AO22X1 U204 ( .IN1(SH[1]), .IN2(n208), .IN3(n210), .IN4(n155), .Q(n174) );
  AO22X1 U205 ( .IN1(SH[1]), .IN2(n207), .IN3(n209), .IN4(n155), .Q(n173) );
  AO22X1 U206 ( .IN1(SH[1]), .IN2(n206), .IN3(n208), .IN4(n155), .Q(n172) );
  AO22X1 U207 ( .IN1(SH[1]), .IN2(n205), .IN3(n207), .IN4(n155), .Q(n171) );
  AO22X1 U208 ( .IN1(SH[1]), .IN2(n204), .IN3(n206), .IN4(n155), .Q(n170) );
  AO22X1 U209 ( .IN1(SH[1]), .IN2(n203), .IN3(n205), .IN4(n155), .Q(n169) );
  AO22X1 U210 ( .IN1(SH[1]), .IN2(n202), .IN3(n204), .IN4(n155), .Q(n168) );
  AO22X1 U211 ( .IN1(SH[1]), .IN2(n201), .IN3(n203), .IN4(n155), .Q(n167) );
  AO22X1 U212 ( .IN1(SH[1]), .IN2(n200), .IN3(n202), .IN4(n155), .Q(n166) );
  AO22X1 U213 ( .IN1(SH[1]), .IN2(n199), .IN3(n201), .IN4(n155), .Q(n165) );
  AO22X1 U214 ( .IN1(SH[1]), .IN2(n198), .IN3(n200), .IN4(n155), .Q(n164) );
  AO22X1 U215 ( .IN1(SH[1]), .IN2(n197), .IN3(n199), .IN4(n155), .Q(n163) );
  AO22X1 U216 ( .IN1(SH[1]), .IN2(n196), .IN3(n198), .IN4(n155), .Q(n162) );
  AO22X1 U217 ( .IN1(SH[1]), .IN2(n195), .IN3(n197), .IN4(n155), .Q(n161) );
  AO22X1 U218 ( .IN1(SH[1]), .IN2(n194), .IN3(n196), .IN4(n155), .Q(n160) );
  AO22X1 U219 ( .IN1(SH[1]), .IN2(n193), .IN3(n195), .IN4(n155), .Q(n159) );
  AND2X1 U220 ( .IN1(n194), .IN2(n155), .Q(n158) );
  AND2X1 U221 ( .IN1(n193), .IN2(n155), .Q(n157) );
  AND2X1 U225 ( .IN1(SH[0]), .IN2(A[31]), .Q(n225) );
  AO22X1 U226 ( .IN1(A[30]), .IN2(SH[0]), .IN3(n191), .IN4(A[31]), .Q(n224) );
  AO22X1 U227 ( .IN1(A[29]), .IN2(SH[0]), .IN3(n191), .IN4(A[30]), .Q(n223) );
  AO22X1 U228 ( .IN1(A[28]), .IN2(SH[0]), .IN3(n191), .IN4(A[29]), .Q(n222) );
  AO22X1 U229 ( .IN1(A[27]), .IN2(SH[0]), .IN3(n191), .IN4(A[28]), .Q(n221) );
  AO22X1 U230 ( .IN1(A[26]), .IN2(SH[0]), .IN3(n191), .IN4(A[27]), .Q(n220) );
  AO22X1 U231 ( .IN1(A[25]), .IN2(SH[0]), .IN3(n191), .IN4(A[26]), .Q(n219) );
  AO22X1 U232 ( .IN1(A[24]), .IN2(SH[0]), .IN3(n191), .IN4(A[25]), .Q(n218) );
  AO22X1 U233 ( .IN1(A[23]), .IN2(SH[0]), .IN3(n191), .IN4(A[24]), .Q(n217) );
  AO22X1 U234 ( .IN1(A[22]), .IN2(SH[0]), .IN3(n191), .IN4(A[23]), .Q(n216) );
  AO22X1 U235 ( .IN1(A[21]), .IN2(SH[0]), .IN3(n191), .IN4(A[22]), .Q(n215) );
  AO22X1 U236 ( .IN1(A[20]), .IN2(SH[0]), .IN3(n191), .IN4(A[21]), .Q(n214) );
  AO22X1 U237 ( .IN1(A[19]), .IN2(SH[0]), .IN3(n191), .IN4(A[20]), .Q(n213) );
  AO22X1 U238 ( .IN1(A[18]), .IN2(SH[0]), .IN3(n191), .IN4(A[19]), .Q(n212) );
  AO22X1 U239 ( .IN1(A[17]), .IN2(SH[0]), .IN3(n191), .IN4(A[18]), .Q(n211) );
  AO22X1 U240 ( .IN1(A[16]), .IN2(SH[0]), .IN3(n191), .IN4(A[17]), .Q(n210) );
  AO22X1 U241 ( .IN1(A[15]), .IN2(SH[0]), .IN3(n191), .IN4(A[16]), .Q(n209) );
  AO22X1 U242 ( .IN1(A[14]), .IN2(SH[0]), .IN3(n191), .IN4(A[15]), .Q(n208) );
  AO22X1 U243 ( .IN1(A[13]), .IN2(SH[0]), .IN3(n191), .IN4(A[14]), .Q(n207) );
  AO22X1 U244 ( .IN1(A[12]), .IN2(SH[0]), .IN3(n191), .IN4(A[13]), .Q(n206) );
  AO22X1 U245 ( .IN1(A[11]), .IN2(SH[0]), .IN3(n191), .IN4(A[12]), .Q(n205) );
  AO22X1 U246 ( .IN1(A[10]), .IN2(SH[0]), .IN3(n191), .IN4(A[11]), .Q(n204) );
  AO22X1 U247 ( .IN1(A[9]), .IN2(SH[0]), .IN3(n191), .IN4(A[10]), .Q(n203) );
  AO22X1 U248 ( .IN1(A[8]), .IN2(SH[0]), .IN3(n191), .IN4(A[9]), .Q(n202) );
  AO22X1 U249 ( .IN1(A[7]), .IN2(SH[0]), .IN3(n191), .IN4(A[8]), .Q(n201) );
  AO22X1 U250 ( .IN1(A[6]), .IN2(SH[0]), .IN3(n191), .IN4(A[7]), .Q(n200) );
  AO22X1 U251 ( .IN1(A[5]), .IN2(SH[0]), .IN3(n191), .IN4(A[6]), .Q(n199) );
  AO22X1 U252 ( .IN1(A[4]), .IN2(SH[0]), .IN3(n191), .IN4(A[5]), .Q(n198) );
  AO22X1 U253 ( .IN1(A[3]), .IN2(SH[0]), .IN3(n191), .IN4(A[4]), .Q(n197) );
  AO22X1 U254 ( .IN1(A[2]), .IN2(SH[0]), .IN3(n191), .IN4(A[3]), .Q(n196) );
  AO22X1 U255 ( .IN1(A[1]), .IN2(SH[0]), .IN3(n191), .IN4(A[2]), .Q(n195) );
  AO22X1 U256 ( .IN1(A[0]), .IN2(SH[0]), .IN3(n191), .IN4(A[1]), .Q(n194) );
  AND2X1 U257 ( .IN1(n191), .IN2(A[0]), .Q(n193) );
  INVX0 U263 ( .INP(SH[1]), .ZN(n155) );
  INVX0 U264 ( .INP(SH[2]), .ZN(n118) );
  INVX0 U265 ( .INP(SH[0]), .ZN(n191) );
  INVX0 U266 ( .INP(SH[3]), .ZN(n81) );
  INVX0 U267 ( .INP(SH[4]), .ZN(n44) );
  INVX0 U268 ( .INP(SH[5]), .ZN(n7) );
  NOR2X0 U269 ( .IN1(SH[7]), .IN2(SH[6]), .QN(n306) );
endmodule


module thumb ( read_instruction_n, instruction_address, instruction, 
        read_data_n, write_data_n, data_address, data, reset_n, clk );
  output [31:0] instruction_address;
  input [15:0] instruction;
  output [31:0] data_address;
  inout [31:0] data;
  input reset_n, clk;
  output read_instruction_n, read_data_n, write_data_n;
  wire   N187, N188, N190, N191, N193, N195, N196, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
         N227, N228, N229, N230, N231, N232, N313, N314, N315, N316, N317,
         N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328,
         N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339,
         N340, N341, N342, N343, N344, \R[7][31] , \R[7][30] , \R[7][29] ,
         \R[7][28] , \R[7][27] , \R[7][26] , \R[7][25] , \R[7][24] ,
         \R[7][23] , \R[7][22] , \R[7][21] , \R[7][20] , \R[7][19] ,
         \R[7][18] , \R[7][17] , \R[7][16] , \R[7][15] , \R[7][14] ,
         \R[7][13] , \R[7][12] , \R[7][11] , \R[7][10] , \R[7][9] , \R[7][8] ,
         \R[7][7] , \R[7][6] , \R[7][5] , \R[7][4] , \R[7][3] , \R[7][2] ,
         \R[7][1] , \R[7][0] , \R[6][31] , \R[6][30] , \R[6][29] , \R[6][28] ,
         \R[6][27] , \R[6][26] , \R[6][25] , \R[6][24] , \R[6][23] ,
         \R[6][22] , \R[6][21] , \R[6][20] , \R[6][19] , \R[6][18] ,
         \R[6][17] , \R[6][16] , \R[6][15] , \R[6][14] , \R[6][13] ,
         \R[6][12] , \R[6][11] , \R[6][10] , \R[6][9] , \R[6][8] , \R[6][7] ,
         \R[6][6] , \R[6][5] , \R[6][4] , \R[6][3] , \R[6][2] , \R[6][1] ,
         \R[6][0] , \R[5][31] , \R[5][30] , \R[5][29] , \R[5][28] , \R[5][27] ,
         \R[5][26] , \R[5][25] , \R[5][24] , \R[5][23] , \R[5][22] ,
         \R[5][21] , \R[5][20] , \R[5][19] , \R[5][18] , \R[5][17] ,
         \R[5][16] , \R[5][15] , \R[5][14] , \R[5][13] , \R[5][12] ,
         \R[5][11] , \R[5][10] , \R[5][9] , \R[5][8] , \R[5][7] , \R[5][6] ,
         \R[5][5] , \R[5][4] , \R[5][3] , \R[5][2] , \R[5][1] , \R[5][0] ,
         \R[4][31] , \R[4][30] , \R[4][29] , \R[4][28] , \R[4][27] ,
         \R[4][26] , \R[4][25] , \R[4][24] , \R[4][23] , \R[4][22] ,
         \R[4][21] , \R[4][20] , \R[4][19] , \R[4][18] , \R[4][17] ,
         \R[4][16] , \R[4][15] , \R[4][14] , \R[4][13] , \R[4][12] ,
         \R[4][11] , \R[4][10] , \R[4][9] , \R[4][8] , \R[4][7] , \R[4][6] ,
         \R[4][5] , \R[4][4] , \R[4][3] , \R[4][2] , \R[4][1] , \R[4][0] ,
         \R[3][31] , \R[3][30] , \R[3][29] , \R[3][28] , \R[3][27] ,
         \R[3][26] , \R[3][25] , \R[3][24] , \R[3][23] , \R[3][22] ,
         \R[3][21] , \R[3][20] , \R[3][19] , \R[3][18] , \R[3][17] ,
         \R[3][16] , \R[3][15] , \R[3][14] , \R[3][13] , \R[3][12] ,
         \R[3][11] , \R[3][10] , \R[3][9] , \R[3][8] , \R[3][7] , \R[3][6] ,
         \R[3][5] , \R[3][4] , \R[3][3] , \R[3][2] , \R[3][1] , \R[3][0] ,
         \R[2][31] , \R[2][30] , \R[2][29] , \R[2][28] , \R[2][27] ,
         \R[2][26] , \R[2][25] , \R[2][24] , \R[2][23] , \R[2][22] ,
         \R[2][21] , \R[2][20] , \R[2][19] , \R[2][18] , \R[2][17] ,
         \R[2][16] , \R[2][15] , \R[2][14] , \R[2][13] , \R[2][12] ,
         \R[2][11] , \R[2][10] , \R[2][9] , \R[2][8] , \R[2][7] , \R[2][6] ,
         \R[2][5] , \R[2][4] , \R[2][3] , \R[2][2] , \R[2][1] , \R[2][0] ,
         \R[1][31] , \R[1][30] , \R[1][29] , \R[1][28] , \R[1][27] ,
         \R[1][26] , \R[1][25] , \R[1][24] , \R[1][23] , \R[1][22] ,
         \R[1][21] , \R[1][20] , \R[1][19] , \R[1][18] , \R[1][17] ,
         \R[1][16] , \R[1][15] , \R[1][14] , \R[1][13] , \R[1][12] ,
         \R[1][11] , \R[1][10] , \R[1][9] , \R[1][8] , \R[1][7] , \R[1][6] ,
         \R[1][5] , \R[1][4] , \R[1][3] , \R[1][2] , \R[1][1] , \R[1][0] ,
         \R[0][31] , \R[0][30] , \R[0][29] , \R[0][28] , \R[0][27] ,
         \R[0][26] , \R[0][25] , \R[0][24] , \R[0][23] , \R[0][22] ,
         \R[0][21] , \R[0][20] , \R[0][19] , \R[0][18] , \R[0][17] ,
         \R[0][16] , \R[0][15] , \R[0][14] , \R[0][13] , \R[0][12] ,
         \R[0][11] , \R[0][10] , \R[0][9] , \R[0][8] , \R[0][7] , \R[0][6] ,
         \R[0][5] , \R[0][4] , \R[0][3] , \R[0][2] , \R[0][1] , \R[0][0] ,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N498, N547, N548, N550,
         N595, N596, N598, N599, N685, N686, N687, N688, N690, N693, N694,
         N695, N767, N768, N769, N771, N772, N773, N777, N1148, N1149, N1150,
         N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160,
         N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170,
         N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180,
         N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192,
         N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202,
         N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212,
         N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222,
         N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232,
         N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242,
         N1243, N1244, N2429, N3556, N3557, N3558, N3559, N3560, N3561, N3562,
         N3563, N3564, N3565, N3566, N3567, N3568, N3569, N3570, N3571, N3572,
         N3573, N3574, N3575, N3576, N3577, N3578, N3579, N3580, N3581, N3582,
         N3583, N3584, N3585, N3586, N3587, N3588, N3654, N3687, N3688, N3689,
         N3690, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3698, N3699,
         N3700, N3701, N3702, N3703, N3704, N3705, N3706, N3707, N3708, N3709,
         N3710, N3711, N3712, N3713, N3714, N3715, N3716, N3717, N3718, N3719,
         N3720, N3724, N3725, N3726, N3727, N3728, N3729, N3730, N3731, N3732,
         N3733, N3734, N3735, N3736, N3737, N3738, N3739, N3740, N3741, N3742,
         N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752,
         N3753, N3754, N3755, N3756, N3790, N3791, N3792, N3793, N3794, N3795,
         N3796, N3797, N3798, N3799, N3800, N3801, N3802, N3803, N3804, N3805,
         N3806, N3807, N3808, N3809, N3810, N3811, N3812, N3813, N3814, N3815,
         N3816, N3817, N3818, N3819, N3820, N3821, N3822, N3826, N3827, N3828,
         N3829, N3830, N3831, N3832, N3833, N3834, N3835, N3836, N3837, N3838,
         N3839, N3840, N3841, N3842, N3843, N3844, N3845, N3846, N3847, N3848,
         N3849, N3850, N3851, N3852, N3853, N3854, N3855, N3856, N3857, N3858,
         N4634, N4637, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, \U3/U74/Z_0 , \U3/U74/Z_1 , \U3/U74/Z_2 , \U3/U74/Z_3 ,
         \U3/U74/Z_4 , \U3/U74/Z_5 , \U3/U74/Z_6 , \U3/U74/Z_7 , \U3/U74/Z_8 ,
         \U3/U74/Z_9 , \U3/U74/Z_10 , \U3/U74/Z_11 , \U3/U74/Z_12 ,
         \U3/U74/Z_13 , \U3/U74/Z_14 , \U3/U74/Z_15 , \U3/U74/Z_16 ,
         \U3/U74/Z_17 , \U3/U74/Z_18 , \U3/U74/Z_19 , \U3/U74/Z_20 ,
         \U3/U74/Z_21 , \U3/U74/Z_22 , \U3/U74/Z_23 , \U3/U74/Z_24 ,
         \U3/U74/Z_25 , \U3/U74/Z_26 , \U3/U74/Z_27 , \U3/U74/Z_28 ,
         \U3/U74/Z_29 , \U3/U74/Z_30 , \U3/U74/Z_31 , \U3/U75/Z_0 ,
         \U3/U75/Z_1 , \U3/U75/Z_2 , \U3/U75/Z_3 , \U3/U75/Z_4 , \U3/U75/Z_5 ,
         \U3/U75/Z_6 , \U3/U75/Z_7 , \U3/U75/Z_8 , \U3/U75/Z_9 , \U3/U75/Z_10 ,
         \U3/U75/Z_11 , \U3/U75/Z_12 , \U3/U75/Z_13 , \U3/U75/Z_14 ,
         \U3/U75/Z_15 , \U3/U75/Z_16 , \U3/U75/Z_17 , \U3/U75/Z_18 ,
         \U3/U75/Z_19 , \U3/U75/Z_20 , \U3/U75/Z_21 , \U3/U75/Z_22 ,
         \U3/U75/Z_23 , \U3/U75/Z_24 , \U3/U75/Z_25 , \U3/U75/Z_26 ,
         \U3/U75/Z_27 , \U3/U75/Z_28 , \U3/U75/Z_29 , \U3/U75/Z_30 ,
         \U3/U75/Z_31 , \U3/U76/Z_0 , \U3/U77/Z_0 , n2988, n2991, n2994, n2995,
         n2996, n3000, n3002, n3004, n3006, n3008, n3010, n3012, n3014, n3016,
         n3018, n3020, n3022, n3024, n3026, n3028, n3030, n3032, n3034, n3036,
         n3038, n3040, n3042, n3044, n3046, n3048, n3050, n3052, n3054, n3056,
         n3058, n3060, n3062, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3096, n3130, n3131, n3132, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3795,
         n3797, n3799, n3800, n3802, \r150/A[3] , n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771;
  wire   [15:0] IF_IR;
  wire   [31:0] IF_PC;
  wire   [7:0] ID_imm_offset;
  wire   [31:0] ID_Rn;
  wire   [31:0] ID_Rd;
  wire   [31:0] ID_Rm_Rs;
  wire   [31:0] ID_PC;
  wire   [31:0] SP;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign read_instruction_n = 1'b0;

  DFFASX1 write_data_n_reg ( .D(N4634), .CLK(clk), .SETB(reset_n), .Q(
        write_data_n), .QN(n5735) );
  DFFASX1 read_data_n_reg ( .D(N4637), .CLK(clk), .SETB(reset_n), .Q(
        read_data_n) );
  DFFX1 \ID_PC_reg[31]  ( .D(IF_PC[31]), .CLK(clk), .Q(ID_PC[31]) );
  DFFARX1 \PC_reg[31]  ( .D(N344), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[31]) );
  DFFX1 \ID_PC_reg[0]  ( .D(IF_PC[0]), .CLK(clk), .Q(ID_PC[0]) );
  DFFARX1 \PC_reg[0]  ( .D(N313), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[0]) );
  DFFX1 \ID_PC_reg[1]  ( .D(IF_PC[1]), .CLK(clk), .Q(ID_PC[1]) );
  DFFARX1 \PC_reg[1]  ( .D(N314), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[1]) );
  DFFX1 \ID_PC_reg[2]  ( .D(IF_PC[2]), .CLK(clk), .Q(ID_PC[2]) );
  DFFARX1 \PC_reg[2]  ( .D(N315), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[2]) );
  DFFX1 \ID_PC_reg[3]  ( .D(IF_PC[3]), .CLK(clk), .Q(ID_PC[3]) );
  DFFARX1 \PC_reg[3]  ( .D(N316), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[3]) );
  DFFX1 \ID_PC_reg[4]  ( .D(IF_PC[4]), .CLK(clk), .Q(ID_PC[4]) );
  DFFARX1 \PC_reg[4]  ( .D(N317), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[4]) );
  DFFX1 \ID_PC_reg[5]  ( .D(IF_PC[5]), .CLK(clk), .Q(ID_PC[5]) );
  DFFARX1 \PC_reg[5]  ( .D(N318), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[5]) );
  DFFX1 \ID_PC_reg[6]  ( .D(IF_PC[6]), .CLK(clk), .Q(ID_PC[6]) );
  DFFARX1 \PC_reg[6]  ( .D(N319), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[6]) );
  DFFX1 \ID_PC_reg[7]  ( .D(IF_PC[7]), .CLK(clk), .Q(ID_PC[7]) );
  DFFARX1 \PC_reg[7]  ( .D(N320), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[7]) );
  DFFX1 \ID_PC_reg[8]  ( .D(IF_PC[8]), .CLK(clk), .Q(ID_PC[8]) );
  DFFARX1 \PC_reg[8]  ( .D(N321), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[8]) );
  DFFX1 \ID_PC_reg[9]  ( .D(IF_PC[9]), .CLK(clk), .Q(ID_PC[9]) );
  DFFARX1 \PC_reg[9]  ( .D(N322), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[9]) );
  DFFX1 \ID_PC_reg[10]  ( .D(IF_PC[10]), .CLK(clk), .Q(ID_PC[10]) );
  DFFARX1 \PC_reg[10]  ( .D(N323), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[10]) );
  DFFX1 \ID_PC_reg[11]  ( .D(IF_PC[11]), .CLK(clk), .Q(ID_PC[11]) );
  DFFARX1 \PC_reg[11]  ( .D(N324), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[11]) );
  DFFX1 \ID_PC_reg[12]  ( .D(IF_PC[12]), .CLK(clk), .Q(ID_PC[12]) );
  DFFARX1 \PC_reg[12]  ( .D(N325), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[12]) );
  DFFX1 \ID_PC_reg[13]  ( .D(IF_PC[13]), .CLK(clk), .Q(ID_PC[13]) );
  DFFARX1 \PC_reg[13]  ( .D(N326), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[13]) );
  DFFX1 \ID_PC_reg[14]  ( .D(IF_PC[14]), .CLK(clk), .Q(ID_PC[14]) );
  DFFARX1 \PC_reg[14]  ( .D(N327), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[14]) );
  DFFX1 \ID_PC_reg[15]  ( .D(IF_PC[15]), .CLK(clk), .Q(ID_PC[15]) );
  DFFARX1 \PC_reg[15]  ( .D(N328), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[15]) );
  DFFX1 \ID_PC_reg[16]  ( .D(IF_PC[16]), .CLK(clk), .Q(ID_PC[16]) );
  DFFARX1 \PC_reg[16]  ( .D(N329), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[16]) );
  DFFX1 \ID_PC_reg[17]  ( .D(IF_PC[17]), .CLK(clk), .Q(ID_PC[17]) );
  DFFARX1 \PC_reg[17]  ( .D(N330), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[17]) );
  DFFX1 \ID_PC_reg[18]  ( .D(IF_PC[18]), .CLK(clk), .Q(ID_PC[18]) );
  DFFARX1 \PC_reg[18]  ( .D(N331), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[18]) );
  DFFX1 \ID_PC_reg[19]  ( .D(IF_PC[19]), .CLK(clk), .Q(ID_PC[19]) );
  DFFARX1 \PC_reg[19]  ( .D(N332), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[19]) );
  DFFX1 \ID_PC_reg[20]  ( .D(IF_PC[20]), .CLK(clk), .Q(ID_PC[20]) );
  DFFARX1 \PC_reg[20]  ( .D(N333), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[20]) );
  DFFX1 \ID_PC_reg[21]  ( .D(IF_PC[21]), .CLK(clk), .Q(ID_PC[21]) );
  DFFARX1 \PC_reg[21]  ( .D(N334), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[21]) );
  DFFX1 \ID_PC_reg[22]  ( .D(IF_PC[22]), .CLK(clk), .Q(ID_PC[22]) );
  DFFARX1 \PC_reg[22]  ( .D(N335), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[22]) );
  DFFX1 \ID_PC_reg[23]  ( .D(IF_PC[23]), .CLK(clk), .Q(ID_PC[23]) );
  DFFARX1 \PC_reg[23]  ( .D(N336), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[23]) );
  DFFX1 \ID_PC_reg[24]  ( .D(IF_PC[24]), .CLK(clk), .Q(ID_PC[24]) );
  DFFARX1 \PC_reg[24]  ( .D(N337), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[24]) );
  DFFX1 \ID_PC_reg[25]  ( .D(IF_PC[25]), .CLK(clk), .Q(ID_PC[25]) );
  DFFARX1 \PC_reg[25]  ( .D(N338), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[25]) );
  DFFX1 \ID_PC_reg[26]  ( .D(IF_PC[26]), .CLK(clk), .Q(ID_PC[26]) );
  DFFARX1 \PC_reg[26]  ( .D(N339), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[26]) );
  DFFX1 \ID_PC_reg[27]  ( .D(IF_PC[27]), .CLK(clk), .Q(ID_PC[27]) );
  DFFARX1 \PC_reg[27]  ( .D(N340), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[27]) );
  DFFX1 \ID_PC_reg[28]  ( .D(IF_PC[28]), .CLK(clk), .Q(ID_PC[28]) );
  DFFARX1 \PC_reg[28]  ( .D(N341), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[28]) );
  DFFX1 \ID_PC_reg[29]  ( .D(IF_PC[29]), .CLK(clk), .Q(ID_PC[29]) );
  DFFARX1 \PC_reg[29]  ( .D(N342), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[29]) );
  DFFX1 \ID_PC_reg[30]  ( .D(IF_PC[30]), .CLK(clk), .Q(ID_PC[30]) );
  DFFARX1 \PC_reg[30]  ( .D(N343), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[30]) );
  DFFARX1 branch_taken_reg ( .D(n3792), .CLK(clk), .RSTB(reset_n), .Q(n3842), 
        .QN(n5711) );
  DFFX1 \IF_IR_reg[9]  ( .D(n3791), .CLK(clk), .Q(N195), .QN(n5727) );
  DFFX1 \IF_IR_reg[10]  ( .D(n3790), .CLK(clk), .Q(N196), .QN(n5726) );
  DFFX1 \IF_IR_reg[11]  ( .D(n3789), .CLK(clk), .Q(IF_IR[11]), .QN(n3799) );
  DFFX1 \IF_IR_reg[12]  ( .D(n3788), .CLK(clk), .Q(IF_IR[12]), .QN(n3797) );
  DFFX1 \IF_IR_reg[14]  ( .D(n3787), .CLK(clk), .Q(IF_IR[14]), .QN(n3132) );
  DFFX1 \IF_IR_reg[15]  ( .D(n3786), .CLK(clk), .Q(IF_IR[15]), .QN(n3131) );
  DFFX1 \IF_IR_reg[13]  ( .D(n3785), .CLK(clk), .Q(IF_IR[13]), .QN(n3130) );
  DFFX1 \ID_Rn_reg[0]  ( .D(n3784), .CLK(clk), .Q(ID_Rn[0]) );
  DFFX1 \ID_Rn_reg[1]  ( .D(n3783), .CLK(clk), .Q(ID_Rn[1]) );
  DFFX1 \ID_Rn_reg[2]  ( .D(n3782), .CLK(clk), .Q(ID_Rn[2]) );
  DFFX1 \ID_Rn_reg[3]  ( .D(n3781), .CLK(clk), .Q(ID_Rn[3]) );
  DFFX1 \ID_Rn_reg[4]  ( .D(n3780), .CLK(clk), .Q(ID_Rn[4]) );
  DFFX1 \ID_Rn_reg[5]  ( .D(n3779), .CLK(clk), .Q(ID_Rn[5]) );
  DFFX1 \ID_Rn_reg[6]  ( .D(n3778), .CLK(clk), .Q(ID_Rn[6]) );
  DFFX1 \ID_Rn_reg[7]  ( .D(n3777), .CLK(clk), .Q(ID_Rn[7]) );
  DFFX1 \ID_Rn_reg[8]  ( .D(n3776), .CLK(clk), .Q(ID_Rn[8]) );
  DFFX1 \ID_Rn_reg[9]  ( .D(n3775), .CLK(clk), .Q(ID_Rn[9]) );
  DFFX1 \ID_Rn_reg[10]  ( .D(n3774), .CLK(clk), .Q(ID_Rn[10]) );
  DFFX1 \ID_Rn_reg[11]  ( .D(n3773), .CLK(clk), .Q(ID_Rn[11]) );
  DFFX1 \ID_Rn_reg[12]  ( .D(n3772), .CLK(clk), .Q(ID_Rn[12]) );
  DFFX1 \ID_Rn_reg[13]  ( .D(n3771), .CLK(clk), .Q(ID_Rn[13]) );
  DFFX1 \ID_Rn_reg[14]  ( .D(n3770), .CLK(clk), .Q(ID_Rn[14]) );
  DFFX1 \ID_Rn_reg[15]  ( .D(n3769), .CLK(clk), .Q(ID_Rn[15]) );
  DFFX1 \ID_Rn_reg[16]  ( .D(n3768), .CLK(clk), .Q(ID_Rn[16]) );
  DFFX1 \ID_Rn_reg[17]  ( .D(n3767), .CLK(clk), .Q(ID_Rn[17]) );
  DFFX1 \ID_Rn_reg[18]  ( .D(n3766), .CLK(clk), .Q(ID_Rn[18]) );
  DFFX1 \ID_Rn_reg[19]  ( .D(n3765), .CLK(clk), .Q(ID_Rn[19]) );
  DFFX1 \ID_Rn_reg[20]  ( .D(n3764), .CLK(clk), .Q(ID_Rn[20]) );
  DFFX1 \ID_Rn_reg[21]  ( .D(n3763), .CLK(clk), .Q(ID_Rn[21]) );
  DFFX1 \ID_Rn_reg[22]  ( .D(n3762), .CLK(clk), .Q(ID_Rn[22]) );
  DFFX1 \ID_Rn_reg[23]  ( .D(n3761), .CLK(clk), .Q(ID_Rn[23]) );
  DFFX1 \ID_Rn_reg[24]  ( .D(n3760), .CLK(clk), .Q(ID_Rn[24]) );
  DFFX1 \ID_Rn_reg[25]  ( .D(n3759), .CLK(clk), .Q(ID_Rn[25]) );
  DFFX1 \ID_Rn_reg[26]  ( .D(n3758), .CLK(clk), .Q(ID_Rn[26]) );
  DFFX1 \ID_Rn_reg[27]  ( .D(n3757), .CLK(clk), .Q(ID_Rn[27]) );
  DFFX1 \ID_Rn_reg[28]  ( .D(n3756), .CLK(clk), .Q(ID_Rn[28]) );
  DFFX1 \ID_Rn_reg[29]  ( .D(n3755), .CLK(clk), .Q(ID_Rn[29]) );
  DFFX1 \ID_Rn_reg[30]  ( .D(n3754), .CLK(clk), .Q(ID_Rn[30]) );
  DFFX1 \ID_Rn_reg[31]  ( .D(n3753), .CLK(clk), .Q(ID_Rn[31]) );
  DFFX1 \ID_opcode_reg[0]  ( .D(n3752), .CLK(clk), .Q(n3803), .QN(\r150/A[3] )
         );
  DFFX1 \ID_opcode_reg[1]  ( .D(n3751), .CLK(clk), .Q(n3843), .QN(n5724) );
  DFFX1 \ID_opcode_reg[2]  ( .D(n3750), .CLK(clk), .Q(n3805), .QN(n5723) );
  DFFX1 \ID_opcode_reg[4]  ( .D(n3749), .CLK(clk), .Q(n3804), .QN(n5722) );
  DFFX1 \EX_opcode_reg[4]  ( .D(n3748), .CLK(clk), .QN(n5706) );
  DFFX1 \ID_opcode_reg[5]  ( .D(n3747), .CLK(clk), .Q(n3844), .QN(n5721) );
  DFFX1 \IF_IR_reg[8]  ( .D(n3746), .CLK(clk), .Q(n5719), .QN(n3800) );
  DFFX1 \IF_IR_reg[7]  ( .D(n3745), .CLK(clk), .Q(N193), .QN(n3096) );
  DFFX1 \ID_imm_offset_reg[7]  ( .D(n3744), .CLK(clk), .Q(ID_imm_offset[7]) );
  DFFX1 \IF_IR_reg[6]  ( .D(n3743), .CLK(clk), .Q(n5705), .QN(n5728) );
  DFFX1 \ID_Rm_Rs_reg[0]  ( .D(n3742), .CLK(clk), .Q(ID_Rm_Rs[0]), .QN(n3094)
         );
  DFFX1 \ID_Rm_Rs_reg[1]  ( .D(n3741), .CLK(clk), .Q(ID_Rm_Rs[1]), .QN(n3093)
         );
  DFFX1 \ID_Rm_Rs_reg[2]  ( .D(n3740), .CLK(clk), .Q(ID_Rm_Rs[2]), .QN(n3092)
         );
  DFFX1 \ID_Rm_Rs_reg[3]  ( .D(n3739), .CLK(clk), .Q(ID_Rm_Rs[3]), .QN(n3091)
         );
  DFFX1 \ID_Rm_Rs_reg[4]  ( .D(n3738), .CLK(clk), .Q(ID_Rm_Rs[4]), .QN(n3090)
         );
  DFFX1 \ID_Rm_Rs_reg[5]  ( .D(n3737), .CLK(clk), .Q(ID_Rm_Rs[5]), .QN(n3089)
         );
  DFFX1 \ID_Rm_Rs_reg[6]  ( .D(n3736), .CLK(clk), .Q(ID_Rm_Rs[6]), .QN(n3088)
         );
  DFFX1 \ID_Rm_Rs_reg[7]  ( .D(n3735), .CLK(clk), .Q(ID_Rm_Rs[7]), .QN(n3087)
         );
  DFFX1 \ID_Rm_Rs_reg[8]  ( .D(n3734), .CLK(clk), .Q(ID_Rm_Rs[8]), .QN(n3086)
         );
  DFFX1 \ID_Rm_Rs_reg[9]  ( .D(n3733), .CLK(clk), .Q(ID_Rm_Rs[9]), .QN(n3085)
         );
  DFFX1 \ID_Rm_Rs_reg[10]  ( .D(n3732), .CLK(clk), .Q(ID_Rm_Rs[10]), .QN(n3084) );
  DFFX1 \ID_Rm_Rs_reg[11]  ( .D(n3731), .CLK(clk), .Q(ID_Rm_Rs[11]), .QN(n3083) );
  DFFX1 \ID_Rm_Rs_reg[12]  ( .D(n3730), .CLK(clk), .Q(ID_Rm_Rs[12]), .QN(n3082) );
  DFFX1 \ID_Rm_Rs_reg[13]  ( .D(n3729), .CLK(clk), .Q(ID_Rm_Rs[13]), .QN(n3081) );
  DFFX1 \ID_Rm_Rs_reg[14]  ( .D(n3728), .CLK(clk), .Q(ID_Rm_Rs[14]), .QN(n3080) );
  DFFX1 \ID_Rm_Rs_reg[15]  ( .D(n3727), .CLK(clk), .Q(ID_Rm_Rs[15]), .QN(n3079) );
  DFFX1 \ID_Rm_Rs_reg[16]  ( .D(n3726), .CLK(clk), .Q(ID_Rm_Rs[16]), .QN(n3078) );
  DFFX1 \ID_Rm_Rs_reg[17]  ( .D(n3725), .CLK(clk), .Q(ID_Rm_Rs[17]), .QN(n3077) );
  DFFX1 \ID_Rm_Rs_reg[18]  ( .D(n3724), .CLK(clk), .Q(ID_Rm_Rs[18]), .QN(n3076) );
  DFFX1 \ID_Rm_Rs_reg[19]  ( .D(n3723), .CLK(clk), .Q(ID_Rm_Rs[19]), .QN(n3075) );
  DFFX1 \ID_Rm_Rs_reg[20]  ( .D(n3722), .CLK(clk), .Q(ID_Rm_Rs[20]), .QN(n3074) );
  DFFX1 \ID_Rm_Rs_reg[21]  ( .D(n3721), .CLK(clk), .Q(ID_Rm_Rs[21]), .QN(n3073) );
  DFFX1 \ID_Rm_Rs_reg[22]  ( .D(n3720), .CLK(clk), .Q(ID_Rm_Rs[22]), .QN(n3072) );
  DFFX1 \ID_Rm_Rs_reg[23]  ( .D(n3719), .CLK(clk), .Q(ID_Rm_Rs[23]), .QN(n3071) );
  DFFX1 \ID_Rm_Rs_reg[24]  ( .D(n3718), .CLK(clk), .Q(ID_Rm_Rs[24]), .QN(n3070) );
  DFFX1 \ID_Rm_Rs_reg[25]  ( .D(n3717), .CLK(clk), .Q(ID_Rm_Rs[25]), .QN(n3069) );
  DFFX1 \ID_Rm_Rs_reg[26]  ( .D(n3716), .CLK(clk), .Q(ID_Rm_Rs[26]), .QN(n3068) );
  DFFX1 \ID_Rm_Rs_reg[27]  ( .D(n3715), .CLK(clk), .Q(ID_Rm_Rs[27]), .QN(n3067) );
  DFFX1 \ID_Rm_Rs_reg[28]  ( .D(n3714), .CLK(clk), .Q(ID_Rm_Rs[28]), .QN(n3066) );
  DFFX1 \ID_Rm_Rs_reg[29]  ( .D(n3713), .CLK(clk), .Q(ID_Rm_Rs[29]), .QN(n3065) );
  DFFX1 \ID_Rm_Rs_reg[30]  ( .D(n3712), .CLK(clk), .Q(ID_Rm_Rs[30]), .QN(n3064) );
  DFFX1 \ID_Rm_Rs_reg[31]  ( .D(n3711), .CLK(clk), .Q(N2429), .QN(n5725) );
  DFFX1 \ID_opcode_reg[3]  ( .D(n3710), .CLK(clk), .Q(n3807), .QN(n5720) );
  DFFX1 \EX_opcode_reg[3]  ( .D(n3709), .CLK(clk), .Q(n3884), .QN(n5710) );
  DFFX1 \ID_Rd_reg[0]  ( .D(n3708), .CLK(clk), .Q(ID_Rd[0]), .QN(n3062) );
  DFFX1 \DR_reg[0]  ( .D(n3707), .CLK(clk), .Q(n5740) );
  DFFX1 \ID_Rd_reg[1]  ( .D(n3706), .CLK(clk), .Q(ID_Rd[1]), .QN(n3060) );
  DFFX1 \DR_reg[1]  ( .D(n3705), .CLK(clk), .Q(n5741) );
  DFFX1 \ID_Rd_reg[2]  ( .D(n3704), .CLK(clk), .Q(ID_Rd[2]), .QN(n3058) );
  DFFX1 \DR_reg[2]  ( .D(n3703), .CLK(clk), .Q(n5742) );
  DFFX1 \ID_Rd_reg[3]  ( .D(n3702), .CLK(clk), .Q(ID_Rd[3]), .QN(n3056) );
  DFFX1 \DR_reg[3]  ( .D(n3701), .CLK(clk), .Q(n5743) );
  DFFX1 \ID_Rd_reg[4]  ( .D(n3700), .CLK(clk), .Q(ID_Rd[4]), .QN(n3054) );
  DFFX1 \DR_reg[4]  ( .D(n3699), .CLK(clk), .Q(n5744) );
  DFFX1 \ID_Rd_reg[5]  ( .D(n3698), .CLK(clk), .Q(ID_Rd[5]), .QN(n3052) );
  DFFX1 \DR_reg[5]  ( .D(n3697), .CLK(clk), .Q(n5745) );
  DFFX1 \ID_Rd_reg[6]  ( .D(n3696), .CLK(clk), .Q(ID_Rd[6]), .QN(n3050) );
  DFFX1 \DR_reg[6]  ( .D(n3695), .CLK(clk), .Q(n5746) );
  DFFX1 \ID_Rd_reg[7]  ( .D(n3694), .CLK(clk), .Q(ID_Rd[7]), .QN(n3048) );
  DFFX1 \DR_reg[7]  ( .D(n3693), .CLK(clk), .Q(n5747) );
  DFFX1 \ID_Rd_reg[8]  ( .D(n3692), .CLK(clk), .Q(ID_Rd[8]), .QN(n3046) );
  DFFX1 \DR_reg[8]  ( .D(n3691), .CLK(clk), .Q(n5748) );
  DFFX1 \ID_Rd_reg[9]  ( .D(n3690), .CLK(clk), .Q(ID_Rd[9]), .QN(n3044) );
  DFFX1 \DR_reg[9]  ( .D(n3689), .CLK(clk), .Q(n5749) );
  DFFX1 \ID_Rd_reg[10]  ( .D(n3688), .CLK(clk), .Q(ID_Rd[10]), .QN(n3042) );
  DFFX1 \DR_reg[10]  ( .D(n3687), .CLK(clk), .Q(n5750) );
  DFFX1 \ID_Rd_reg[11]  ( .D(n3686), .CLK(clk), .Q(ID_Rd[11]), .QN(n3040) );
  DFFX1 \DR_reg[11]  ( .D(n3685), .CLK(clk), .Q(n5751) );
  DFFX1 \ID_Rd_reg[12]  ( .D(n3684), .CLK(clk), .Q(ID_Rd[12]), .QN(n3038) );
  DFFX1 \DR_reg[12]  ( .D(n3683), .CLK(clk), .Q(n5752) );
  DFFX1 \ID_Rd_reg[13]  ( .D(n3682), .CLK(clk), .Q(ID_Rd[13]), .QN(n3036) );
  DFFX1 \DR_reg[13]  ( .D(n3681), .CLK(clk), .Q(n5753) );
  DFFX1 \ID_Rd_reg[14]  ( .D(n3680), .CLK(clk), .Q(ID_Rd[14]), .QN(n3034) );
  DFFX1 \DR_reg[14]  ( .D(n3679), .CLK(clk), .Q(n5754) );
  DFFX1 \ID_Rd_reg[15]  ( .D(n3678), .CLK(clk), .Q(ID_Rd[15]), .QN(n3032) );
  DFFX1 \DR_reg[15]  ( .D(n3677), .CLK(clk), .Q(n5755) );
  DFFX1 \ID_Rd_reg[16]  ( .D(n3676), .CLK(clk), .Q(ID_Rd[16]), .QN(n3030) );
  DFFX1 \DR_reg[16]  ( .D(n3675), .CLK(clk), .Q(n5756) );
  DFFX1 \ID_Rd_reg[17]  ( .D(n3674), .CLK(clk), .Q(ID_Rd[17]), .QN(n3028) );
  DFFX1 \DR_reg[17]  ( .D(n3673), .CLK(clk), .Q(n5757) );
  DFFX1 \ID_Rd_reg[18]  ( .D(n3672), .CLK(clk), .Q(ID_Rd[18]), .QN(n3026) );
  DFFX1 \DR_reg[18]  ( .D(n3671), .CLK(clk), .Q(n5758) );
  DFFX1 \ID_Rd_reg[19]  ( .D(n3670), .CLK(clk), .Q(ID_Rd[19]), .QN(n3024) );
  DFFX1 \DR_reg[19]  ( .D(n3669), .CLK(clk), .Q(n5759) );
  DFFX1 \ID_Rd_reg[20]  ( .D(n3668), .CLK(clk), .Q(ID_Rd[20]), .QN(n3022) );
  DFFX1 \DR_reg[20]  ( .D(n3667), .CLK(clk), .Q(n5760) );
  DFFX1 \ID_Rd_reg[21]  ( .D(n3666), .CLK(clk), .Q(ID_Rd[21]), .QN(n3020) );
  DFFX1 \DR_reg[21]  ( .D(n3665), .CLK(clk), .Q(n5761) );
  DFFX1 \ID_Rd_reg[22]  ( .D(n3664), .CLK(clk), .Q(ID_Rd[22]), .QN(n3018) );
  DFFX1 \DR_reg[22]  ( .D(n3663), .CLK(clk), .Q(n5762) );
  DFFX1 \ID_Rd_reg[23]  ( .D(n3662), .CLK(clk), .Q(ID_Rd[23]), .QN(n3016) );
  DFFX1 \DR_reg[23]  ( .D(n3661), .CLK(clk), .Q(n5763) );
  DFFX1 \ID_Rd_reg[24]  ( .D(n3660), .CLK(clk), .Q(ID_Rd[24]), .QN(n3014) );
  DFFX1 \DR_reg[24]  ( .D(n3659), .CLK(clk), .Q(n5764) );
  DFFX1 \ID_Rd_reg[25]  ( .D(n3658), .CLK(clk), .Q(ID_Rd[25]), .QN(n3012) );
  DFFX1 \DR_reg[25]  ( .D(n3657), .CLK(clk), .Q(n5765) );
  DFFX1 \ID_Rd_reg[26]  ( .D(n3656), .CLK(clk), .Q(ID_Rd[26]), .QN(n3010) );
  DFFX1 \DR_reg[26]  ( .D(n3655), .CLK(clk), .Q(n5766) );
  DFFX1 \ID_Rd_reg[27]  ( .D(n3654), .CLK(clk), .Q(ID_Rd[27]), .QN(n3008) );
  DFFX1 \DR_reg[27]  ( .D(n3653), .CLK(clk), .Q(n5767) );
  DFFX1 \ID_Rd_reg[28]  ( .D(n3652), .CLK(clk), .Q(ID_Rd[28]), .QN(n3006) );
  DFFX1 \DR_reg[28]  ( .D(n3651), .CLK(clk), .Q(n5768) );
  DFFX1 \ID_Rd_reg[29]  ( .D(n3650), .CLK(clk), .Q(ID_Rd[29]), .QN(n3004) );
  DFFX1 \DR_reg[29]  ( .D(n3649), .CLK(clk), .Q(n5769) );
  DFFX1 \ID_Rd_reg[30]  ( .D(n3648), .CLK(clk), .Q(ID_Rd[30]), .QN(n3002) );
  DFFX1 \DR_reg[30]  ( .D(n3647), .CLK(clk), .Q(n5770) );
  DFFX1 \ID_Rd_reg[31]  ( .D(n3646), .CLK(clk), .Q(ID_Rd[31]), .QN(n3000) );
  DFFX1 \DR_reg[31]  ( .D(n3645), .CLK(clk), .Q(n5771) );
  DFFX1 \ID_imm_offset_reg[6]  ( .D(n3644), .CLK(clk), .Q(ID_imm_offset[6]) );
  DFFX1 \IF_IR_reg[5]  ( .D(n3643), .CLK(clk), .Q(N188), .QN(n5732) );
  DFFX1 \ID_imm_offset_reg[5]  ( .D(n3642), .CLK(clk), .Q(ID_imm_offset[5]) );
  DFFX1 \IF_IR_reg[4]  ( .D(n3641), .CLK(clk), .Q(N187), .QN(n5733) );
  DFFX1 \ID_imm_offset_reg[4]  ( .D(n3640), .CLK(clk), .Q(ID_imm_offset[4]), 
        .QN(n2996) );
  DFFX1 \IF_IR_reg[3]  ( .D(n3639), .CLK(clk), .Q(n5718), .QN(n5734) );
  DFFX1 \IF_IR_reg[2]  ( .D(n3637), .CLK(clk), .Q(N191), .QN(n5729) );
  DFFX1 \ID_Rd_code_reg[2]  ( .D(n3635), .CLK(clk), .Q(n3880) );
  DFFX1 \EX_Rd_code_reg[2]  ( .D(n3634), .CLK(clk), .Q(n3808), .QN(n5717) );
  DFFX1 \IF_IR_reg[1]  ( .D(n3633), .CLK(clk), .Q(N190), .QN(n5730) );
  DFFX1 \ID_Rd_code_reg[1]  ( .D(n3631), .CLK(clk), .Q(n3881) );
  DFFX1 \EX_Rd_code_reg[1]  ( .D(n3630), .CLK(clk), .Q(n3806), .QN(n5716) );
  DFFX1 \IF_IR_reg[0]  ( .D(n3629), .CLK(clk), .Q(n5715), .QN(n5731) );
  DFFX1 \ID_Rd_code_reg[0]  ( .D(n3627), .CLK(clk), .Q(n3809) );
  DFFX1 \EX_Rd_code_reg[0]  ( .D(n3626), .CLK(clk), .Q(n3883), .QN(n5714) );
  DFFX1 \EX_opcode_reg[5]  ( .D(n3625), .CLK(clk), .Q(n3845), .QN(n5709) );
  DFFX1 \EX_opcode_reg[2]  ( .D(n3624), .CLK(clk), .Q(n3846), .QN(n5707) );
  DFFX1 \EX_opcode_reg[1]  ( .D(n3623), .CLK(clk), .Q(n3882), .QN(n5708) );
  DFFX1 \EX_opcode_reg[0]  ( .D(n3622), .CLK(clk), .QN(n5713) );
  DFFX1 C_Flag_reg ( .D(n3621), .CLK(clk), .Q(n3917), .QN(n5712) );
  DFFX1 \branch_target_reg[0]  ( .D(n3620), .CLK(clk), .Q(n3879) );
  DFFX1 \branch_target_reg[1]  ( .D(n3619), .CLK(clk), .Q(n3878) );
  DFFX1 \branch_target_reg[2]  ( .D(n3618), .CLK(clk), .Q(n3877) );
  DFFX1 \branch_target_reg[3]  ( .D(n3617), .CLK(clk), .Q(n3876) );
  DFFX1 \branch_target_reg[4]  ( .D(n3616), .CLK(clk), .Q(n3875) );
  DFFX1 \branch_target_reg[5]  ( .D(n3615), .CLK(clk), .Q(n3874) );
  DFFX1 \branch_target_reg[6]  ( .D(n3614), .CLK(clk), .Q(n3873) );
  DFFX1 \branch_target_reg[7]  ( .D(n3613), .CLK(clk), .Q(n3872) );
  DFFX1 \branch_target_reg[8]  ( .D(n3612), .CLK(clk), .Q(n3871) );
  DFFX1 \branch_target_reg[9]  ( .D(n3611), .CLK(clk), .Q(n3870) );
  DFFX1 \branch_target_reg[10]  ( .D(n3610), .CLK(clk), .Q(n3869) );
  DFFX1 \branch_target_reg[11]  ( .D(n3609), .CLK(clk), .Q(n3868) );
  DFFX1 \branch_target_reg[12]  ( .D(n3608), .CLK(clk), .Q(n3867) );
  DFFX1 \branch_target_reg[13]  ( .D(n3607), .CLK(clk), .Q(n3866) );
  DFFX1 \branch_target_reg[14]  ( .D(n3606), .CLK(clk), .Q(n3865) );
  DFFX1 \branch_target_reg[15]  ( .D(n3605), .CLK(clk), .Q(n3864) );
  DFFX1 \branch_target_reg[16]  ( .D(n3604), .CLK(clk), .Q(n3863) );
  DFFX1 \branch_target_reg[17]  ( .D(n3603), .CLK(clk), .Q(n3862) );
  DFFX1 \branch_target_reg[18]  ( .D(n3602), .CLK(clk), .Q(n3861) );
  DFFX1 \branch_target_reg[19]  ( .D(n3601), .CLK(clk), .Q(n3860) );
  DFFX1 \branch_target_reg[20]  ( .D(n3600), .CLK(clk), .Q(n3859) );
  DFFX1 \branch_target_reg[21]  ( .D(n3599), .CLK(clk), .Q(n3858) );
  DFFX1 \branch_target_reg[22]  ( .D(n3598), .CLK(clk), .Q(n3857) );
  DFFX1 \branch_target_reg[23]  ( .D(n3597), .CLK(clk), .Q(n3856) );
  DFFX1 \branch_target_reg[24]  ( .D(n3596), .CLK(clk), .Q(n3855) );
  DFFX1 \branch_target_reg[25]  ( .D(n3595), .CLK(clk), .Q(n3854) );
  DFFX1 \branch_target_reg[26]  ( .D(n3594), .CLK(clk), .Q(n3853) );
  DFFX1 \branch_target_reg[27]  ( .D(n3593), .CLK(clk), .Q(n3852) );
  DFFX1 \branch_target_reg[28]  ( .D(n3592), .CLK(clk), .Q(n3851) );
  DFFX1 \branch_target_reg[29]  ( .D(n3591), .CLK(clk), .Q(n3850) );
  DFFX1 \branch_target_reg[30]  ( .D(n3590), .CLK(clk), .Q(n3849) );
  DFFX1 \branch_target_reg[31]  ( .D(n3589), .CLK(clk), .Q(n3848) );
  DFFX1 \IF_PC_reg[31]  ( .D(n3588), .CLK(clk), .Q(IF_PC[31]) );
  DFFX1 \IF_PC_reg[0]  ( .D(n3587), .CLK(clk), .Q(IF_PC[0]) );
  DFFX1 \IF_PC_reg[1]  ( .D(n3586), .CLK(clk), .Q(IF_PC[1]) );
  DFFX1 \IF_PC_reg[2]  ( .D(n3585), .CLK(clk), .Q(IF_PC[2]) );
  DFFX1 \IF_PC_reg[3]  ( .D(n3584), .CLK(clk), .Q(IF_PC[3]) );
  DFFX1 \IF_PC_reg[4]  ( .D(n3583), .CLK(clk), .Q(IF_PC[4]) );
  DFFX1 \IF_PC_reg[5]  ( .D(n3582), .CLK(clk), .Q(IF_PC[5]) );
  DFFX1 \IF_PC_reg[6]  ( .D(n3581), .CLK(clk), .Q(IF_PC[6]) );
  DFFX1 \IF_PC_reg[7]  ( .D(n3580), .CLK(clk), .Q(IF_PC[7]) );
  DFFX1 \IF_PC_reg[8]  ( .D(n3579), .CLK(clk), .Q(IF_PC[8]) );
  DFFX1 \IF_PC_reg[9]  ( .D(n3578), .CLK(clk), .Q(IF_PC[9]) );
  DFFX1 \IF_PC_reg[10]  ( .D(n3577), .CLK(clk), .Q(IF_PC[10]) );
  DFFX1 \IF_PC_reg[11]  ( .D(n3576), .CLK(clk), .Q(IF_PC[11]) );
  DFFX1 \IF_PC_reg[12]  ( .D(n3575), .CLK(clk), .Q(IF_PC[12]) );
  DFFX1 \IF_PC_reg[13]  ( .D(n3574), .CLK(clk), .Q(IF_PC[13]) );
  DFFX1 \IF_PC_reg[14]  ( .D(n3573), .CLK(clk), .Q(IF_PC[14]) );
  DFFX1 \IF_PC_reg[15]  ( .D(n3572), .CLK(clk), .Q(IF_PC[15]) );
  DFFX1 \IF_PC_reg[16]  ( .D(n3571), .CLK(clk), .Q(IF_PC[16]) );
  DFFX1 \IF_PC_reg[17]  ( .D(n3570), .CLK(clk), .Q(IF_PC[17]) );
  DFFX1 \IF_PC_reg[18]  ( .D(n3569), .CLK(clk), .Q(IF_PC[18]) );
  DFFX1 \IF_PC_reg[19]  ( .D(n3568), .CLK(clk), .Q(IF_PC[19]) );
  DFFX1 \IF_PC_reg[20]  ( .D(n3567), .CLK(clk), .Q(IF_PC[20]) );
  DFFX1 \IF_PC_reg[21]  ( .D(n3566), .CLK(clk), .Q(IF_PC[21]) );
  DFFX1 \IF_PC_reg[22]  ( .D(n3565), .CLK(clk), .Q(IF_PC[22]) );
  DFFX1 \IF_PC_reg[23]  ( .D(n3564), .CLK(clk), .Q(IF_PC[23]) );
  DFFX1 \IF_PC_reg[24]  ( .D(n3563), .CLK(clk), .Q(IF_PC[24]) );
  DFFX1 \IF_PC_reg[25]  ( .D(n3562), .CLK(clk), .Q(IF_PC[25]) );
  DFFX1 \IF_PC_reg[26]  ( .D(n3561), .CLK(clk), .Q(IF_PC[26]) );
  DFFX1 \IF_PC_reg[27]  ( .D(n3560), .CLK(clk), .Q(IF_PC[27]) );
  DFFX1 \IF_PC_reg[28]  ( .D(n3559), .CLK(clk), .Q(IF_PC[28]) );
  DFFX1 \IF_PC_reg[29]  ( .D(n3558), .CLK(clk), .Q(IF_PC[29]) );
  DFFX1 \IF_PC_reg[30]  ( .D(n3557), .CLK(clk), .Q(IF_PC[30]) );
  DFFX1 \SP_reg[31]  ( .D(n3556), .CLK(clk), .Q(SP[31]) );
  DFFX1 \ALU_out_reg[0]  ( .D(n3555), .CLK(clk), .Q(n3810) );
  DFFX1 \data_address_reg[0]  ( .D(n3554), .CLK(clk), .Q(data_address[0]) );
  DFFX1 \SP_reg[0]  ( .D(n3553), .CLK(clk), .Q(SP[0]) );
  DFFX1 \EX_ALU_out_reg[0]  ( .D(n3552), .CLK(clk), .Q(n3916) );
  DFFX1 \ALU_out_reg[1]  ( .D(n3551), .CLK(clk), .Q(n3811) );
  DFFX1 \data_address_reg[1]  ( .D(n3550), .CLK(clk), .Q(data_address[1]) );
  DFFX1 \SP_reg[1]  ( .D(n3549), .CLK(clk), .Q(SP[1]) );
  DFFX1 \EX_ALU_out_reg[1]  ( .D(n3548), .CLK(clk), .Q(n3915) );
  DFFX1 \ALU_out_reg[2]  ( .D(n3547), .CLK(clk), .Q(n3812) );
  DFFX1 \data_address_reg[2]  ( .D(n3546), .CLK(clk), .Q(data_address[2]) );
  DFFX1 \SP_reg[2]  ( .D(n3545), .CLK(clk), .Q(SP[2]) );
  DFFX1 \EX_ALU_out_reg[2]  ( .D(n3544), .CLK(clk), .Q(n3914) );
  DFFX1 \ALU_out_reg[3]  ( .D(n3543), .CLK(clk), .Q(n3813) );
  DFFX1 \data_address_reg[3]  ( .D(n3542), .CLK(clk), .Q(data_address[3]) );
  DFFX1 \SP_reg[3]  ( .D(n3541), .CLK(clk), .Q(SP[3]) );
  DFFX1 \EX_ALU_out_reg[3]  ( .D(n3540), .CLK(clk), .Q(n3913) );
  DFFX1 \ALU_out_reg[4]  ( .D(n3539), .CLK(clk), .Q(n3814) );
  DFFX1 \data_address_reg[4]  ( .D(n3538), .CLK(clk), .Q(data_address[4]) );
  DFFX1 \SP_reg[4]  ( .D(n3537), .CLK(clk), .Q(SP[4]) );
  DFFX1 \EX_ALU_out_reg[4]  ( .D(n3536), .CLK(clk), .Q(n3912) );
  DFFX1 \ALU_out_reg[5]  ( .D(n3535), .CLK(clk), .Q(n3815) );
  DFFX1 \data_address_reg[5]  ( .D(n3534), .CLK(clk), .Q(data_address[5]) );
  DFFX1 \SP_reg[5]  ( .D(n3533), .CLK(clk), .Q(SP[5]) );
  DFFX1 \EX_ALU_out_reg[5]  ( .D(n3532), .CLK(clk), .Q(n3911) );
  DFFX1 \ALU_out_reg[6]  ( .D(n3531), .CLK(clk), .Q(n3816) );
  DFFX1 \data_address_reg[6]  ( .D(n3530), .CLK(clk), .Q(data_address[6]) );
  DFFX1 \SP_reg[6]  ( .D(n3529), .CLK(clk), .Q(SP[6]) );
  DFFX1 \EX_ALU_out_reg[6]  ( .D(n3528), .CLK(clk), .Q(n3910) );
  DFFX1 \ALU_out_reg[7]  ( .D(n3527), .CLK(clk), .Q(n3817) );
  DFFX1 \data_address_reg[7]  ( .D(n3526), .CLK(clk), .Q(data_address[7]) );
  DFFX1 \SP_reg[7]  ( .D(n3525), .CLK(clk), .Q(SP[7]) );
  DFFX1 \EX_ALU_out_reg[7]  ( .D(n3524), .CLK(clk), .Q(n3909) );
  DFFX1 \ALU_out_reg[8]  ( .D(n3523), .CLK(clk), .Q(n3818) );
  DFFX1 \data_address_reg[8]  ( .D(n3522), .CLK(clk), .Q(data_address[8]) );
  DFFX1 \SP_reg[8]  ( .D(n3521), .CLK(clk), .Q(SP[8]) );
  DFFX1 \EX_ALU_out_reg[8]  ( .D(n3520), .CLK(clk), .Q(n3908) );
  DFFX1 \ALU_out_reg[9]  ( .D(n3519), .CLK(clk), .Q(n3819) );
  DFFX1 \data_address_reg[9]  ( .D(n3518), .CLK(clk), .Q(data_address[9]) );
  DFFX1 \SP_reg[9]  ( .D(n3517), .CLK(clk), .Q(SP[9]) );
  DFFX1 \EX_ALU_out_reg[9]  ( .D(n3516), .CLK(clk), .Q(n3907) );
  DFFX1 \ALU_out_reg[10]  ( .D(n3515), .CLK(clk), .Q(n3820) );
  DFFX1 \data_address_reg[10]  ( .D(n3514), .CLK(clk), .Q(data_address[10]) );
  DFFX1 \SP_reg[10]  ( .D(n3513), .CLK(clk), .Q(SP[10]) );
  DFFX1 \EX_ALU_out_reg[10]  ( .D(n3512), .CLK(clk), .Q(n3906) );
  DFFX1 \ALU_out_reg[11]  ( .D(n3511), .CLK(clk), .Q(n3821) );
  DFFX1 \data_address_reg[11]  ( .D(n3510), .CLK(clk), .Q(data_address[11]) );
  DFFX1 \SP_reg[11]  ( .D(n3509), .CLK(clk), .Q(SP[11]) );
  DFFX1 \EX_ALU_out_reg[11]  ( .D(n3508), .CLK(clk), .Q(n3905) );
  DFFX1 \ALU_out_reg[12]  ( .D(n3507), .CLK(clk), .Q(n3822) );
  DFFX1 \data_address_reg[12]  ( .D(n3506), .CLK(clk), .Q(data_address[12]) );
  DFFX1 \SP_reg[12]  ( .D(n3505), .CLK(clk), .Q(SP[12]) );
  DFFX1 \EX_ALU_out_reg[12]  ( .D(n3504), .CLK(clk), .Q(n3904) );
  DFFX1 \ALU_out_reg[13]  ( .D(n3503), .CLK(clk), .Q(n3823) );
  DFFX1 \data_address_reg[13]  ( .D(n3502), .CLK(clk), .Q(data_address[13]) );
  DFFX1 \SP_reg[13]  ( .D(n3501), .CLK(clk), .Q(SP[13]) );
  DFFX1 \EX_ALU_out_reg[13]  ( .D(n3500), .CLK(clk), .Q(n3903) );
  DFFX1 \ALU_out_reg[14]  ( .D(n3499), .CLK(clk), .Q(n3824) );
  DFFX1 \data_address_reg[14]  ( .D(n3498), .CLK(clk), .Q(data_address[14]) );
  DFFX1 \SP_reg[14]  ( .D(n3497), .CLK(clk), .Q(SP[14]) );
  DFFX1 \EX_ALU_out_reg[14]  ( .D(n3496), .CLK(clk), .Q(n3902) );
  DFFX1 \ALU_out_reg[15]  ( .D(n3495), .CLK(clk), .Q(n3825) );
  DFFX1 \data_address_reg[15]  ( .D(n3494), .CLK(clk), .Q(data_address[15]) );
  DFFX1 \SP_reg[15]  ( .D(n3493), .CLK(clk), .Q(SP[15]) );
  DFFX1 \EX_ALU_out_reg[15]  ( .D(n3492), .CLK(clk), .Q(n3901) );
  DFFX1 \ALU_out_reg[16]  ( .D(n3491), .CLK(clk), .Q(n3826) );
  DFFX1 \data_address_reg[16]  ( .D(n3490), .CLK(clk), .Q(data_address[16]) );
  DFFX1 \SP_reg[16]  ( .D(n3489), .CLK(clk), .Q(SP[16]) );
  DFFX1 \EX_ALU_out_reg[16]  ( .D(n3488), .CLK(clk), .Q(n3900) );
  DFFX1 \ALU_out_reg[17]  ( .D(n3487), .CLK(clk), .Q(n3827) );
  DFFX1 \data_address_reg[17]  ( .D(n3486), .CLK(clk), .Q(data_address[17]) );
  DFFX1 \SP_reg[17]  ( .D(n3485), .CLK(clk), .Q(SP[17]) );
  DFFX1 \EX_ALU_out_reg[17]  ( .D(n3484), .CLK(clk), .Q(n3899) );
  DFFX1 \ALU_out_reg[18]  ( .D(n3483), .CLK(clk), .Q(n3828) );
  DFFX1 \data_address_reg[18]  ( .D(n3482), .CLK(clk), .Q(data_address[18]) );
  DFFX1 \SP_reg[18]  ( .D(n3481), .CLK(clk), .Q(SP[18]) );
  DFFX1 \EX_ALU_out_reg[18]  ( .D(n3480), .CLK(clk), .Q(n3898) );
  DFFX1 \ALU_out_reg[19]  ( .D(n3479), .CLK(clk), .Q(n3829) );
  DFFX1 \data_address_reg[19]  ( .D(n3478), .CLK(clk), .Q(data_address[19]) );
  DFFX1 \SP_reg[19]  ( .D(n3477), .CLK(clk), .Q(SP[19]) );
  DFFX1 \EX_ALU_out_reg[19]  ( .D(n3476), .CLK(clk), .Q(n3897) );
  DFFX1 \ALU_out_reg[20]  ( .D(n3475), .CLK(clk), .Q(n3830) );
  DFFX1 \data_address_reg[20]  ( .D(n3474), .CLK(clk), .Q(data_address[20]) );
  DFFX1 \SP_reg[20]  ( .D(n3473), .CLK(clk), .Q(SP[20]) );
  DFFX1 \EX_ALU_out_reg[20]  ( .D(n3472), .CLK(clk), .Q(n3896) );
  DFFX1 \ALU_out_reg[21]  ( .D(n3471), .CLK(clk), .Q(n3831) );
  DFFX1 \data_address_reg[21]  ( .D(n3470), .CLK(clk), .Q(data_address[21]) );
  DFFX1 \SP_reg[21]  ( .D(n3469), .CLK(clk), .Q(SP[21]) );
  DFFX1 \EX_ALU_out_reg[21]  ( .D(n3468), .CLK(clk), .Q(n3895) );
  DFFX1 \ALU_out_reg[22]  ( .D(n3467), .CLK(clk), .Q(n3832) );
  DFFX1 \data_address_reg[22]  ( .D(n3466), .CLK(clk), .Q(data_address[22]) );
  DFFX1 \SP_reg[22]  ( .D(n3465), .CLK(clk), .Q(SP[22]) );
  DFFX1 \EX_ALU_out_reg[22]  ( .D(n3464), .CLK(clk), .Q(n3894) );
  DFFX1 \ALU_out_reg[23]  ( .D(n3463), .CLK(clk), .Q(n3833) );
  DFFX1 \data_address_reg[23]  ( .D(n3462), .CLK(clk), .Q(data_address[23]) );
  DFFX1 \SP_reg[23]  ( .D(n3461), .CLK(clk), .Q(SP[23]) );
  DFFX1 \EX_ALU_out_reg[23]  ( .D(n3460), .CLK(clk), .Q(n3893) );
  DFFX1 \ALU_out_reg[24]  ( .D(n3459), .CLK(clk), .Q(n3834) );
  DFFX1 \data_address_reg[24]  ( .D(n3458), .CLK(clk), .Q(data_address[24]) );
  DFFX1 \SP_reg[24]  ( .D(n3457), .CLK(clk), .Q(SP[24]) );
  DFFX1 \EX_ALU_out_reg[24]  ( .D(n3456), .CLK(clk), .Q(n3892) );
  DFFX1 \ALU_out_reg[25]  ( .D(n3455), .CLK(clk), .Q(n3835) );
  DFFX1 \data_address_reg[25]  ( .D(n3454), .CLK(clk), .Q(data_address[25]) );
  DFFX1 \SP_reg[25]  ( .D(n3453), .CLK(clk), .Q(SP[25]) );
  DFFX1 \EX_ALU_out_reg[25]  ( .D(n3452), .CLK(clk), .Q(n3891) );
  DFFX1 \ALU_out_reg[26]  ( .D(n3451), .CLK(clk), .Q(n3836) );
  DFFX1 \data_address_reg[26]  ( .D(n3450), .CLK(clk), .Q(data_address[26]) );
  DFFX1 \SP_reg[26]  ( .D(n3449), .CLK(clk), .Q(SP[26]) );
  DFFX1 \EX_ALU_out_reg[26]  ( .D(n3448), .CLK(clk), .Q(n3890) );
  DFFX1 \ALU_out_reg[27]  ( .D(n3447), .CLK(clk), .Q(n3837) );
  DFFX1 \data_address_reg[27]  ( .D(n3446), .CLK(clk), .Q(data_address[27]) );
  DFFX1 \SP_reg[27]  ( .D(n3445), .CLK(clk), .Q(SP[27]) );
  DFFX1 \EX_ALU_out_reg[27]  ( .D(n3444), .CLK(clk), .Q(n3889) );
  DFFX1 \ALU_out_reg[28]  ( .D(n3443), .CLK(clk), .Q(n3838) );
  DFFX1 \data_address_reg[28]  ( .D(n3442), .CLK(clk), .Q(data_address[28]) );
  DFFX1 \SP_reg[28]  ( .D(n3441), .CLK(clk), .Q(SP[28]) );
  DFFX1 \EX_ALU_out_reg[28]  ( .D(n3440), .CLK(clk), .Q(n3888) );
  DFFX1 \ALU_out_reg[29]  ( .D(n3439), .CLK(clk), .Q(n3839) );
  DFFX1 \data_address_reg[29]  ( .D(n3438), .CLK(clk), .Q(data_address[29]) );
  DFFX1 \SP_reg[29]  ( .D(n3437), .CLK(clk), .Q(SP[29]) );
  DFFX1 \EX_ALU_out_reg[29]  ( .D(n3436), .CLK(clk), .Q(n3887) );
  DFFX1 \ALU_out_reg[30]  ( .D(n3435), .CLK(clk), .Q(n3840) );
  DFFX1 \data_address_reg[30]  ( .D(n3434), .CLK(clk), .Q(data_address[30]) );
  DFFX1 \SP_reg[30]  ( .D(n3433), .CLK(clk), .Q(SP[30]) );
  DFFX1 \EX_ALU_out_reg[30]  ( .D(n3432), .CLK(clk), .Q(n3886) );
  DFFX1 \ALU_out_reg[31]  ( .D(n3431), .CLK(clk), .Q(n3841) );
  DFFX1 \data_address_reg[31]  ( .D(n3430), .CLK(clk), .Q(data_address[31]) );
  DFFX1 \EX_ALU_out_reg[31]  ( .D(n3429), .CLK(clk), .Q(n3885) );
  DFFX1 \ALU_out_reg[32]  ( .D(n3428), .CLK(clk), .Q(n3847) );
  DFFASX1 \R_reg[7][31]  ( .D(n3427), .CLK(clk), .SETB(reset_n), .Q(\R[7][31] ) );
  DFFASX1 \R_reg[7][30]  ( .D(n3426), .CLK(clk), .SETB(reset_n), .Q(\R[7][30] ) );
  DFFASX1 \R_reg[7][29]  ( .D(n3425), .CLK(clk), .SETB(reset_n), .Q(\R[7][29] ) );
  DFFASX1 \R_reg[7][28]  ( .D(n3424), .CLK(clk), .SETB(reset_n), .Q(\R[7][28] ) );
  DFFASX1 \R_reg[7][27]  ( .D(n3423), .CLK(clk), .SETB(reset_n), .Q(\R[7][27] ) );
  DFFASX1 \R_reg[7][26]  ( .D(n3422), .CLK(clk), .SETB(reset_n), .Q(\R[7][26] ) );
  DFFASX1 \R_reg[7][25]  ( .D(n3421), .CLK(clk), .SETB(reset_n), .Q(\R[7][25] ) );
  DFFASX1 \R_reg[7][24]  ( .D(n3420), .CLK(clk), .SETB(reset_n), .Q(\R[7][24] ) );
  DFFASX1 \R_reg[7][23]  ( .D(n3419), .CLK(clk), .SETB(reset_n), .Q(\R[7][23] ) );
  DFFASX1 \R_reg[7][22]  ( .D(n3418), .CLK(clk), .SETB(reset_n), .Q(\R[7][22] ) );
  DFFASX1 \R_reg[7][21]  ( .D(n3417), .CLK(clk), .SETB(reset_n), .Q(\R[7][21] ) );
  DFFASX1 \R_reg[7][20]  ( .D(n3416), .CLK(clk), .SETB(reset_n), .Q(\R[7][20] ) );
  DFFASX1 \R_reg[7][19]  ( .D(n3415), .CLK(clk), .SETB(reset_n), .Q(\R[7][19] ) );
  DFFASX1 \R_reg[7][18]  ( .D(n3414), .CLK(clk), .SETB(reset_n), .Q(\R[7][18] ) );
  DFFASX1 \R_reg[7][17]  ( .D(n3413), .CLK(clk), .SETB(reset_n), .Q(\R[7][17] ) );
  DFFASX1 \R_reg[7][16]  ( .D(n3412), .CLK(clk), .SETB(reset_n), .Q(\R[7][16] ) );
  DFFASX1 \R_reg[7][15]  ( .D(n3411), .CLK(clk), .SETB(reset_n), .Q(\R[7][15] ) );
  DFFASX1 \R_reg[7][14]  ( .D(n3410), .CLK(clk), .SETB(reset_n), .Q(\R[7][14] ) );
  DFFASX1 \R_reg[7][13]  ( .D(n3409), .CLK(clk), .SETB(reset_n), .Q(\R[7][13] ) );
  DFFASX1 \R_reg[7][12]  ( .D(n3408), .CLK(clk), .SETB(reset_n), .Q(\R[7][12] ) );
  DFFASX1 \R_reg[7][11]  ( .D(n3407), .CLK(clk), .SETB(reset_n), .Q(\R[7][11] ) );
  DFFASX1 \R_reg[7][10]  ( .D(n3406), .CLK(clk), .SETB(reset_n), .Q(\R[7][10] ) );
  DFFASX1 \R_reg[7][9]  ( .D(n3405), .CLK(clk), .SETB(reset_n), .Q(\R[7][9] )
         );
  DFFASX1 \R_reg[7][8]  ( .D(n3404), .CLK(clk), .SETB(reset_n), .Q(\R[7][8] )
         );
  DFFASX1 \R_reg[7][7]  ( .D(n3403), .CLK(clk), .SETB(reset_n), .Q(\R[7][7] )
         );
  DFFASX1 \R_reg[7][6]  ( .D(n3402), .CLK(clk), .SETB(reset_n), .Q(\R[7][6] )
         );
  DFFASX1 \R_reg[7][5]  ( .D(n3401), .CLK(clk), .SETB(reset_n), .Q(\R[7][5] )
         );
  DFFASX1 \R_reg[7][4]  ( .D(n3400), .CLK(clk), .SETB(reset_n), .Q(\R[7][4] )
         );
  DFFASX1 \R_reg[7][3]  ( .D(n3399), .CLK(clk), .SETB(reset_n), .Q(\R[7][3] )
         );
  DFFASX1 \R_reg[7][2]  ( .D(n3398), .CLK(clk), .SETB(reset_n), .Q(\R[7][2] )
         );
  DFFASX1 \R_reg[7][1]  ( .D(n3397), .CLK(clk), .SETB(reset_n), .Q(\R[7][1] )
         );
  DFFASX1 \R_reg[7][0]  ( .D(n3396), .CLK(clk), .SETB(reset_n), .Q(\R[7][0] )
         );
  DFFASX1 \R_reg[6][31]  ( .D(n3395), .CLK(clk), .SETB(reset_n), .Q(\R[6][31] ) );
  DFFASX1 \R_reg[6][30]  ( .D(n3394), .CLK(clk), .SETB(reset_n), .Q(\R[6][30] ) );
  DFFASX1 \R_reg[6][29]  ( .D(n3393), .CLK(clk), .SETB(reset_n), .Q(\R[6][29] ) );
  DFFASX1 \R_reg[6][28]  ( .D(n3392), .CLK(clk), .SETB(reset_n), .Q(\R[6][28] ) );
  DFFASX1 \R_reg[6][27]  ( .D(n3391), .CLK(clk), .SETB(reset_n), .Q(\R[6][27] ) );
  DFFASX1 \R_reg[6][26]  ( .D(n3390), .CLK(clk), .SETB(reset_n), .Q(\R[6][26] ) );
  DFFASX1 \R_reg[6][25]  ( .D(n3389), .CLK(clk), .SETB(reset_n), .Q(\R[6][25] ) );
  DFFASX1 \R_reg[6][24]  ( .D(n3388), .CLK(clk), .SETB(reset_n), .Q(\R[6][24] ) );
  DFFASX1 \R_reg[6][23]  ( .D(n3387), .CLK(clk), .SETB(reset_n), .Q(\R[6][23] ) );
  DFFASX1 \R_reg[6][22]  ( .D(n3386), .CLK(clk), .SETB(reset_n), .Q(\R[6][22] ) );
  DFFASX1 \R_reg[6][21]  ( .D(n3385), .CLK(clk), .SETB(reset_n), .Q(\R[6][21] ) );
  DFFASX1 \R_reg[6][20]  ( .D(n3384), .CLK(clk), .SETB(reset_n), .Q(\R[6][20] ) );
  DFFASX1 \R_reg[6][19]  ( .D(n3383), .CLK(clk), .SETB(reset_n), .Q(\R[6][19] ) );
  DFFASX1 \R_reg[6][18]  ( .D(n3382), .CLK(clk), .SETB(reset_n), .Q(\R[6][18] ) );
  DFFASX1 \R_reg[6][17]  ( .D(n3381), .CLK(clk), .SETB(reset_n), .Q(\R[6][17] ) );
  DFFASX1 \R_reg[6][16]  ( .D(n3380), .CLK(clk), .SETB(reset_n), .Q(\R[6][16] ) );
  DFFASX1 \R_reg[6][15]  ( .D(n3379), .CLK(clk), .SETB(reset_n), .Q(\R[6][15] ) );
  DFFASX1 \R_reg[6][14]  ( .D(n3378), .CLK(clk), .SETB(reset_n), .Q(\R[6][14] ) );
  DFFASX1 \R_reg[6][13]  ( .D(n3377), .CLK(clk), .SETB(reset_n), .Q(\R[6][13] ) );
  DFFASX1 \R_reg[6][12]  ( .D(n3376), .CLK(clk), .SETB(reset_n), .Q(\R[6][12] ) );
  DFFASX1 \R_reg[6][11]  ( .D(n3375), .CLK(clk), .SETB(reset_n), .Q(\R[6][11] ) );
  DFFASX1 \R_reg[6][10]  ( .D(n3374), .CLK(clk), .SETB(reset_n), .Q(\R[6][10] ) );
  DFFASX1 \R_reg[6][9]  ( .D(n3373), .CLK(clk), .SETB(reset_n), .Q(\R[6][9] )
         );
  DFFASX1 \R_reg[6][8]  ( .D(n3372), .CLK(clk), .SETB(reset_n), .Q(\R[6][8] )
         );
  DFFASX1 \R_reg[6][7]  ( .D(n3371), .CLK(clk), .SETB(reset_n), .Q(\R[6][7] )
         );
  DFFASX1 \R_reg[6][6]  ( .D(n3370), .CLK(clk), .SETB(reset_n), .Q(\R[6][6] )
         );
  DFFASX1 \R_reg[6][5]  ( .D(n3369), .CLK(clk), .SETB(reset_n), .Q(\R[6][5] )
         );
  DFFASX1 \R_reg[6][4]  ( .D(n3368), .CLK(clk), .SETB(reset_n), .Q(\R[6][4] )
         );
  DFFASX1 \R_reg[6][3]  ( .D(n3367), .CLK(clk), .SETB(reset_n), .Q(\R[6][3] )
         );
  DFFASX1 \R_reg[6][2]  ( .D(n3366), .CLK(clk), .SETB(reset_n), .Q(\R[6][2] )
         );
  DFFASX1 \R_reg[6][1]  ( .D(n3365), .CLK(clk), .SETB(reset_n), .Q(\R[6][1] )
         );
  DFFASX1 \R_reg[6][0]  ( .D(n3364), .CLK(clk), .SETB(reset_n), .Q(\R[6][0] )
         );
  DFFASX1 \R_reg[5][31]  ( .D(n3363), .CLK(clk), .SETB(reset_n), .Q(\R[5][31] ) );
  DFFASX1 \R_reg[5][30]  ( .D(n3362), .CLK(clk), .SETB(reset_n), .Q(\R[5][30] ) );
  DFFASX1 \R_reg[5][29]  ( .D(n3361), .CLK(clk), .SETB(reset_n), .Q(\R[5][29] ) );
  DFFASX1 \R_reg[5][28]  ( .D(n3360), .CLK(clk), .SETB(reset_n), .Q(\R[5][28] ) );
  DFFASX1 \R_reg[5][27]  ( .D(n3359), .CLK(clk), .SETB(reset_n), .Q(\R[5][27] ) );
  DFFASX1 \R_reg[5][26]  ( .D(n3358), .CLK(clk), .SETB(reset_n), .Q(\R[5][26] ) );
  DFFASX1 \R_reg[5][25]  ( .D(n3357), .CLK(clk), .SETB(reset_n), .Q(\R[5][25] ) );
  DFFASX1 \R_reg[5][24]  ( .D(n3356), .CLK(clk), .SETB(reset_n), .Q(\R[5][24] ) );
  DFFASX1 \R_reg[5][23]  ( .D(n3355), .CLK(clk), .SETB(reset_n), .Q(\R[5][23] ) );
  DFFASX1 \R_reg[5][22]  ( .D(n3354), .CLK(clk), .SETB(reset_n), .Q(\R[5][22] ) );
  DFFASX1 \R_reg[5][21]  ( .D(n3353), .CLK(clk), .SETB(reset_n), .Q(\R[5][21] ) );
  DFFASX1 \R_reg[5][20]  ( .D(n3352), .CLK(clk), .SETB(reset_n), .Q(\R[5][20] ) );
  DFFASX1 \R_reg[5][19]  ( .D(n3351), .CLK(clk), .SETB(reset_n), .Q(\R[5][19] ) );
  DFFASX1 \R_reg[5][18]  ( .D(n3350), .CLK(clk), .SETB(reset_n), .Q(\R[5][18] ) );
  DFFASX1 \R_reg[5][17]  ( .D(n3349), .CLK(clk), .SETB(reset_n), .Q(\R[5][17] ) );
  DFFASX1 \R_reg[5][16]  ( .D(n3348), .CLK(clk), .SETB(reset_n), .Q(\R[5][16] ) );
  DFFASX1 \R_reg[5][15]  ( .D(n3347), .CLK(clk), .SETB(reset_n), .Q(\R[5][15] ) );
  DFFASX1 \R_reg[5][14]  ( .D(n3346), .CLK(clk), .SETB(reset_n), .Q(\R[5][14] ) );
  DFFASX1 \R_reg[5][13]  ( .D(n3345), .CLK(clk), .SETB(reset_n), .Q(\R[5][13] ) );
  DFFASX1 \R_reg[5][12]  ( .D(n3344), .CLK(clk), .SETB(reset_n), .Q(\R[5][12] ) );
  DFFASX1 \R_reg[5][11]  ( .D(n3343), .CLK(clk), .SETB(reset_n), .Q(\R[5][11] ) );
  DFFASX1 \R_reg[5][10]  ( .D(n3342), .CLK(clk), .SETB(reset_n), .Q(\R[5][10] ) );
  DFFASX1 \R_reg[5][9]  ( .D(n3341), .CLK(clk), .SETB(reset_n), .Q(\R[5][9] )
         );
  DFFASX1 \R_reg[5][8]  ( .D(n3340), .CLK(clk), .SETB(reset_n), .Q(\R[5][8] )
         );
  DFFASX1 \R_reg[5][7]  ( .D(n3339), .CLK(clk), .SETB(reset_n), .Q(\R[5][7] )
         );
  DFFASX1 \R_reg[5][6]  ( .D(n3338), .CLK(clk), .SETB(reset_n), .Q(\R[5][6] )
         );
  DFFASX1 \R_reg[5][5]  ( .D(n3337), .CLK(clk), .SETB(reset_n), .Q(\R[5][5] )
         );
  DFFASX1 \R_reg[5][4]  ( .D(n3336), .CLK(clk), .SETB(reset_n), .Q(\R[5][4] )
         );
  DFFASX1 \R_reg[5][3]  ( .D(n3335), .CLK(clk), .SETB(reset_n), .Q(\R[5][3] )
         );
  DFFASX1 \R_reg[5][2]  ( .D(n3334), .CLK(clk), .SETB(reset_n), .Q(\R[5][2] )
         );
  DFFASX1 \R_reg[5][1]  ( .D(n3333), .CLK(clk), .SETB(reset_n), .Q(\R[5][1] )
         );
  DFFASX1 \R_reg[5][0]  ( .D(n3332), .CLK(clk), .SETB(reset_n), .Q(\R[5][0] )
         );
  DFFASX1 \R_reg[4][31]  ( .D(n3331), .CLK(clk), .SETB(reset_n), .Q(\R[4][31] ) );
  DFFASX1 \R_reg[4][30]  ( .D(n3330), .CLK(clk), .SETB(reset_n), .Q(\R[4][30] ) );
  DFFASX1 \R_reg[4][29]  ( .D(n3329), .CLK(clk), .SETB(reset_n), .Q(\R[4][29] ) );
  DFFASX1 \R_reg[4][28]  ( .D(n3328), .CLK(clk), .SETB(reset_n), .Q(\R[4][28] ) );
  DFFASX1 \R_reg[4][27]  ( .D(n3327), .CLK(clk), .SETB(reset_n), .Q(\R[4][27] ) );
  DFFASX1 \R_reg[4][26]  ( .D(n3326), .CLK(clk), .SETB(reset_n), .Q(\R[4][26] ) );
  DFFASX1 \R_reg[4][25]  ( .D(n3325), .CLK(clk), .SETB(reset_n), .Q(\R[4][25] ) );
  DFFASX1 \R_reg[4][24]  ( .D(n3324), .CLK(clk), .SETB(reset_n), .Q(\R[4][24] ) );
  DFFASX1 \R_reg[4][23]  ( .D(n3323), .CLK(clk), .SETB(reset_n), .Q(\R[4][23] ) );
  DFFASX1 \R_reg[4][22]  ( .D(n3322), .CLK(clk), .SETB(reset_n), .Q(\R[4][22] ) );
  DFFASX1 \R_reg[4][21]  ( .D(n3321), .CLK(clk), .SETB(reset_n), .Q(\R[4][21] ) );
  DFFASX1 \R_reg[4][20]  ( .D(n3320), .CLK(clk), .SETB(reset_n), .Q(\R[4][20] ) );
  DFFASX1 \R_reg[4][19]  ( .D(n3319), .CLK(clk), .SETB(reset_n), .Q(\R[4][19] ) );
  DFFASX1 \R_reg[4][18]  ( .D(n3318), .CLK(clk), .SETB(reset_n), .Q(\R[4][18] ) );
  DFFASX1 \R_reg[4][17]  ( .D(n3317), .CLK(clk), .SETB(reset_n), .Q(\R[4][17] ) );
  DFFASX1 \R_reg[4][16]  ( .D(n3316), .CLK(clk), .SETB(reset_n), .Q(\R[4][16] ) );
  DFFASX1 \R_reg[4][15]  ( .D(n3315), .CLK(clk), .SETB(reset_n), .Q(\R[4][15] ) );
  DFFASX1 \R_reg[4][14]  ( .D(n3314), .CLK(clk), .SETB(reset_n), .Q(\R[4][14] ) );
  DFFASX1 \R_reg[4][13]  ( .D(n3313), .CLK(clk), .SETB(reset_n), .Q(\R[4][13] ) );
  DFFASX1 \R_reg[4][12]  ( .D(n3312), .CLK(clk), .SETB(reset_n), .Q(\R[4][12] ) );
  DFFASX1 \R_reg[4][11]  ( .D(n3311), .CLK(clk), .SETB(reset_n), .Q(\R[4][11] ) );
  DFFASX1 \R_reg[4][10]  ( .D(n3310), .CLK(clk), .SETB(reset_n), .Q(\R[4][10] ) );
  DFFASX1 \R_reg[4][9]  ( .D(n3309), .CLK(clk), .SETB(reset_n), .Q(\R[4][9] )
         );
  DFFASX1 \R_reg[4][8]  ( .D(n3308), .CLK(clk), .SETB(reset_n), .Q(\R[4][8] )
         );
  DFFASX1 \R_reg[4][7]  ( .D(n3307), .CLK(clk), .SETB(reset_n), .Q(\R[4][7] )
         );
  DFFASX1 \R_reg[4][6]  ( .D(n3306), .CLK(clk), .SETB(reset_n), .Q(\R[4][6] )
         );
  DFFASX1 \R_reg[4][5]  ( .D(n3305), .CLK(clk), .SETB(reset_n), .Q(\R[4][5] )
         );
  DFFASX1 \R_reg[4][4]  ( .D(n3304), .CLK(clk), .SETB(reset_n), .Q(\R[4][4] )
         );
  DFFASX1 \R_reg[4][3]  ( .D(n3303), .CLK(clk), .SETB(reset_n), .Q(\R[4][3] )
         );
  DFFASX1 \R_reg[4][2]  ( .D(n3302), .CLK(clk), .SETB(reset_n), .Q(\R[4][2] )
         );
  DFFASX1 \R_reg[4][1]  ( .D(n3301), .CLK(clk), .SETB(reset_n), .Q(\R[4][1] )
         );
  DFFASX1 \R_reg[4][0]  ( .D(n3300), .CLK(clk), .SETB(reset_n), .Q(\R[4][0] )
         );
  DFFASX1 \R_reg[3][31]  ( .D(n3299), .CLK(clk), .SETB(reset_n), .Q(\R[3][31] ) );
  DFFASX1 \R_reg[3][30]  ( .D(n3298), .CLK(clk), .SETB(reset_n), .Q(\R[3][30] ) );
  DFFASX1 \R_reg[3][29]  ( .D(n3297), .CLK(clk), .SETB(reset_n), .Q(\R[3][29] ) );
  DFFASX1 \R_reg[3][28]  ( .D(n3296), .CLK(clk), .SETB(reset_n), .Q(\R[3][28] ) );
  DFFASX1 \R_reg[3][27]  ( .D(n3295), .CLK(clk), .SETB(reset_n), .Q(\R[3][27] ) );
  DFFASX1 \R_reg[3][26]  ( .D(n3294), .CLK(clk), .SETB(reset_n), .Q(\R[3][26] ) );
  DFFASX1 \R_reg[3][25]  ( .D(n3293), .CLK(clk), .SETB(reset_n), .Q(\R[3][25] ) );
  DFFASX1 \R_reg[3][24]  ( .D(n3292), .CLK(clk), .SETB(reset_n), .Q(\R[3][24] ) );
  DFFASX1 \R_reg[3][23]  ( .D(n3291), .CLK(clk), .SETB(reset_n), .Q(\R[3][23] ) );
  DFFASX1 \R_reg[3][22]  ( .D(n3290), .CLK(clk), .SETB(reset_n), .Q(\R[3][22] ) );
  DFFASX1 \R_reg[3][21]  ( .D(n3289), .CLK(clk), .SETB(reset_n), .Q(\R[3][21] ) );
  DFFASX1 \R_reg[3][20]  ( .D(n3288), .CLK(clk), .SETB(reset_n), .Q(\R[3][20] ) );
  DFFASX1 \R_reg[3][19]  ( .D(n3287), .CLK(clk), .SETB(reset_n), .Q(\R[3][19] ) );
  DFFASX1 \R_reg[3][18]  ( .D(n3286), .CLK(clk), .SETB(reset_n), .Q(\R[3][18] ) );
  DFFASX1 \R_reg[3][17]  ( .D(n3285), .CLK(clk), .SETB(reset_n), .Q(\R[3][17] ) );
  DFFASX1 \R_reg[3][16]  ( .D(n3284), .CLK(clk), .SETB(reset_n), .Q(\R[3][16] ) );
  DFFASX1 \R_reg[3][15]  ( .D(n3283), .CLK(clk), .SETB(reset_n), .Q(\R[3][15] ) );
  DFFASX1 \R_reg[3][14]  ( .D(n3282), .CLK(clk), .SETB(reset_n), .Q(\R[3][14] ) );
  DFFASX1 \R_reg[3][13]  ( .D(n3281), .CLK(clk), .SETB(reset_n), .Q(\R[3][13] ) );
  DFFASX1 \R_reg[3][12]  ( .D(n3280), .CLK(clk), .SETB(reset_n), .Q(\R[3][12] ) );
  DFFASX1 \R_reg[3][11]  ( .D(n3279), .CLK(clk), .SETB(reset_n), .Q(\R[3][11] ) );
  DFFASX1 \R_reg[3][10]  ( .D(n3278), .CLK(clk), .SETB(reset_n), .Q(\R[3][10] ) );
  DFFASX1 \R_reg[3][9]  ( .D(n3277), .CLK(clk), .SETB(reset_n), .Q(\R[3][9] )
         );
  DFFASX1 \R_reg[3][8]  ( .D(n3276), .CLK(clk), .SETB(reset_n), .Q(\R[3][8] )
         );
  DFFASX1 \R_reg[3][7]  ( .D(n3275), .CLK(clk), .SETB(reset_n), .Q(\R[3][7] )
         );
  DFFASX1 \R_reg[3][6]  ( .D(n3274), .CLK(clk), .SETB(reset_n), .Q(\R[3][6] )
         );
  DFFASX1 \R_reg[3][5]  ( .D(n3273), .CLK(clk), .SETB(reset_n), .Q(\R[3][5] )
         );
  DFFASX1 \R_reg[3][4]  ( .D(n3272), .CLK(clk), .SETB(reset_n), .Q(\R[3][4] )
         );
  DFFASX1 \R_reg[3][3]  ( .D(n3271), .CLK(clk), .SETB(reset_n), .Q(\R[3][3] )
         );
  DFFASX1 \R_reg[3][2]  ( .D(n3270), .CLK(clk), .SETB(reset_n), .Q(\R[3][2] )
         );
  DFFASX1 \R_reg[3][1]  ( .D(n3269), .CLK(clk), .SETB(reset_n), .Q(\R[3][1] )
         );
  DFFASX1 \R_reg[3][0]  ( .D(n3268), .CLK(clk), .SETB(reset_n), .Q(\R[3][0] )
         );
  DFFASX1 \R_reg[2][31]  ( .D(n3267), .CLK(clk), .SETB(reset_n), .Q(\R[2][31] ) );
  DFFASX1 \R_reg[2][30]  ( .D(n3266), .CLK(clk), .SETB(reset_n), .Q(\R[2][30] ) );
  DFFASX1 \R_reg[2][29]  ( .D(n3265), .CLK(clk), .SETB(reset_n), .Q(\R[2][29] ) );
  DFFASX1 \R_reg[2][28]  ( .D(n3264), .CLK(clk), .SETB(reset_n), .Q(\R[2][28] ) );
  DFFASX1 \R_reg[2][27]  ( .D(n3263), .CLK(clk), .SETB(reset_n), .Q(\R[2][27] ) );
  DFFASX1 \R_reg[2][26]  ( .D(n3262), .CLK(clk), .SETB(reset_n), .Q(\R[2][26] ) );
  DFFASX1 \R_reg[2][25]  ( .D(n3261), .CLK(clk), .SETB(reset_n), .Q(\R[2][25] ) );
  DFFASX1 \R_reg[2][24]  ( .D(n3260), .CLK(clk), .SETB(reset_n), .Q(\R[2][24] ) );
  DFFASX1 \R_reg[2][23]  ( .D(n3259), .CLK(clk), .SETB(reset_n), .Q(\R[2][23] ) );
  DFFASX1 \R_reg[2][22]  ( .D(n3258), .CLK(clk), .SETB(reset_n), .Q(\R[2][22] ) );
  DFFASX1 \R_reg[2][21]  ( .D(n3257), .CLK(clk), .SETB(reset_n), .Q(\R[2][21] ) );
  DFFASX1 \R_reg[2][20]  ( .D(n3256), .CLK(clk), .SETB(reset_n), .Q(\R[2][20] ) );
  DFFASX1 \R_reg[2][19]  ( .D(n3255), .CLK(clk), .SETB(reset_n), .Q(\R[2][19] ) );
  DFFASX1 \R_reg[2][18]  ( .D(n3254), .CLK(clk), .SETB(reset_n), .Q(\R[2][18] ) );
  DFFASX1 \R_reg[2][17]  ( .D(n3253), .CLK(clk), .SETB(reset_n), .Q(\R[2][17] ) );
  DFFASX1 \R_reg[2][16]  ( .D(n3252), .CLK(clk), .SETB(reset_n), .Q(\R[2][16] ) );
  DFFASX1 \R_reg[2][15]  ( .D(n3251), .CLK(clk), .SETB(reset_n), .Q(\R[2][15] ) );
  DFFASX1 \R_reg[2][14]  ( .D(n3250), .CLK(clk), .SETB(reset_n), .Q(\R[2][14] ) );
  DFFASX1 \R_reg[2][13]  ( .D(n3249), .CLK(clk), .SETB(reset_n), .Q(\R[2][13] ) );
  DFFASX1 \R_reg[2][12]  ( .D(n3248), .CLK(clk), .SETB(reset_n), .Q(\R[2][12] ) );
  DFFASX1 \R_reg[2][11]  ( .D(n3247), .CLK(clk), .SETB(reset_n), .Q(\R[2][11] ) );
  DFFASX1 \R_reg[2][10]  ( .D(n3246), .CLK(clk), .SETB(reset_n), .Q(\R[2][10] ) );
  DFFASX1 \R_reg[2][9]  ( .D(n3245), .CLK(clk), .SETB(reset_n), .Q(\R[2][9] )
         );
  DFFASX1 \R_reg[2][8]  ( .D(n3244), .CLK(clk), .SETB(reset_n), .Q(\R[2][8] )
         );
  DFFASX1 \R_reg[2][7]  ( .D(n3243), .CLK(clk), .SETB(reset_n), .Q(\R[2][7] )
         );
  DFFASX1 \R_reg[2][6]  ( .D(n3242), .CLK(clk), .SETB(reset_n), .Q(\R[2][6] )
         );
  DFFASX1 \R_reg[2][5]  ( .D(n3241), .CLK(clk), .SETB(reset_n), .Q(\R[2][5] )
         );
  DFFASX1 \R_reg[2][4]  ( .D(n3240), .CLK(clk), .SETB(reset_n), .Q(\R[2][4] )
         );
  DFFASX1 \R_reg[2][3]  ( .D(n3239), .CLK(clk), .SETB(reset_n), .Q(\R[2][3] )
         );
  DFFASX1 \R_reg[2][2]  ( .D(n3238), .CLK(clk), .SETB(reset_n), .Q(\R[2][2] )
         );
  DFFASX1 \R_reg[2][1]  ( .D(n3237), .CLK(clk), .SETB(reset_n), .Q(\R[2][1] )
         );
  DFFASX1 \R_reg[2][0]  ( .D(n3236), .CLK(clk), .SETB(reset_n), .Q(\R[2][0] )
         );
  DFFASX1 \R_reg[1][31]  ( .D(n3235), .CLK(clk), .SETB(reset_n), .Q(\R[1][31] ) );
  DFFASX1 \R_reg[1][30]  ( .D(n3234), .CLK(clk), .SETB(reset_n), .Q(\R[1][30] ) );
  DFFASX1 \R_reg[1][29]  ( .D(n3233), .CLK(clk), .SETB(reset_n), .Q(\R[1][29] ) );
  DFFASX1 \R_reg[1][28]  ( .D(n3232), .CLK(clk), .SETB(reset_n), .Q(\R[1][28] ) );
  DFFASX1 \R_reg[1][27]  ( .D(n3231), .CLK(clk), .SETB(reset_n), .Q(\R[1][27] ) );
  DFFASX1 \R_reg[1][26]  ( .D(n3230), .CLK(clk), .SETB(reset_n), .Q(\R[1][26] ) );
  DFFASX1 \R_reg[1][25]  ( .D(n3229), .CLK(clk), .SETB(reset_n), .Q(\R[1][25] ) );
  DFFASX1 \R_reg[1][24]  ( .D(n3228), .CLK(clk), .SETB(reset_n), .Q(\R[1][24] ) );
  DFFASX1 \R_reg[1][23]  ( .D(n3227), .CLK(clk), .SETB(reset_n), .Q(\R[1][23] ) );
  DFFASX1 \R_reg[1][22]  ( .D(n3226), .CLK(clk), .SETB(reset_n), .Q(\R[1][22] ) );
  DFFASX1 \R_reg[1][21]  ( .D(n3225), .CLK(clk), .SETB(reset_n), .Q(\R[1][21] ) );
  DFFASX1 \R_reg[1][20]  ( .D(n3224), .CLK(clk), .SETB(reset_n), .Q(\R[1][20] ) );
  DFFASX1 \R_reg[1][19]  ( .D(n3223), .CLK(clk), .SETB(reset_n), .Q(\R[1][19] ) );
  DFFASX1 \R_reg[1][18]  ( .D(n3222), .CLK(clk), .SETB(reset_n), .Q(\R[1][18] ) );
  DFFASX1 \R_reg[1][17]  ( .D(n3221), .CLK(clk), .SETB(reset_n), .Q(\R[1][17] ) );
  DFFASX1 \R_reg[1][16]  ( .D(n3220), .CLK(clk), .SETB(reset_n), .Q(\R[1][16] ) );
  DFFASX1 \R_reg[1][15]  ( .D(n3219), .CLK(clk), .SETB(reset_n), .Q(\R[1][15] ) );
  DFFASX1 \R_reg[1][14]  ( .D(n3218), .CLK(clk), .SETB(reset_n), .Q(\R[1][14] ) );
  DFFASX1 \R_reg[1][13]  ( .D(n3217), .CLK(clk), .SETB(reset_n), .Q(\R[1][13] ) );
  DFFASX1 \R_reg[1][12]  ( .D(n3216), .CLK(clk), .SETB(reset_n), .Q(\R[1][12] ) );
  DFFASX1 \R_reg[1][11]  ( .D(n3215), .CLK(clk), .SETB(reset_n), .Q(\R[1][11] ) );
  DFFASX1 \R_reg[1][10]  ( .D(n3214), .CLK(clk), .SETB(reset_n), .Q(\R[1][10] ) );
  DFFASX1 \R_reg[1][9]  ( .D(n3213), .CLK(clk), .SETB(reset_n), .Q(\R[1][9] )
         );
  DFFASX1 \R_reg[1][8]  ( .D(n3212), .CLK(clk), .SETB(reset_n), .Q(\R[1][8] )
         );
  DFFASX1 \R_reg[1][7]  ( .D(n3211), .CLK(clk), .SETB(reset_n), .Q(\R[1][7] )
         );
  DFFASX1 \R_reg[1][6]  ( .D(n3210), .CLK(clk), .SETB(reset_n), .Q(\R[1][6] )
         );
  DFFASX1 \R_reg[1][5]  ( .D(n3209), .CLK(clk), .SETB(reset_n), .Q(\R[1][5] )
         );
  DFFASX1 \R_reg[1][4]  ( .D(n3208), .CLK(clk), .SETB(reset_n), .Q(\R[1][4] )
         );
  DFFASX1 \R_reg[1][3]  ( .D(n3207), .CLK(clk), .SETB(reset_n), .Q(\R[1][3] )
         );
  DFFASX1 \R_reg[1][2]  ( .D(n3206), .CLK(clk), .SETB(reset_n), .Q(\R[1][2] )
         );
  DFFASX1 \R_reg[1][1]  ( .D(n3205), .CLK(clk), .SETB(reset_n), .Q(\R[1][1] )
         );
  DFFASX1 \R_reg[1][0]  ( .D(n3204), .CLK(clk), .SETB(reset_n), .Q(\R[1][0] )
         );
  DFFASX1 \R_reg[0][31]  ( .D(n3203), .CLK(clk), .SETB(reset_n), .Q(\R[0][31] ) );
  DFFASX1 \R_reg[0][30]  ( .D(n3202), .CLK(clk), .SETB(reset_n), .Q(\R[0][30] ) );
  DFFASX1 \R_reg[0][29]  ( .D(n3201), .CLK(clk), .SETB(reset_n), .Q(\R[0][29] ) );
  DFFASX1 \R_reg[0][28]  ( .D(n3200), .CLK(clk), .SETB(reset_n), .Q(\R[0][28] ) );
  DFFASX1 \R_reg[0][27]  ( .D(n3199), .CLK(clk), .SETB(reset_n), .Q(\R[0][27] ) );
  DFFASX1 \R_reg[0][26]  ( .D(n3198), .CLK(clk), .SETB(reset_n), .Q(\R[0][26] ) );
  DFFASX1 \R_reg[0][25]  ( .D(n3197), .CLK(clk), .SETB(reset_n), .Q(\R[0][25] ) );
  DFFASX1 \R_reg[0][24]  ( .D(n3196), .CLK(clk), .SETB(reset_n), .Q(\R[0][24] ) );
  DFFASX1 \R_reg[0][23]  ( .D(n3195), .CLK(clk), .SETB(reset_n), .Q(\R[0][23] ) );
  DFFASX1 \R_reg[0][22]  ( .D(n3194), .CLK(clk), .SETB(reset_n), .Q(\R[0][22] ) );
  DFFASX1 \R_reg[0][21]  ( .D(n3193), .CLK(clk), .SETB(reset_n), .Q(\R[0][21] ) );
  DFFASX1 \R_reg[0][20]  ( .D(n3192), .CLK(clk), .SETB(reset_n), .Q(\R[0][20] ) );
  DFFASX1 \R_reg[0][19]  ( .D(n3191), .CLK(clk), .SETB(reset_n), .Q(\R[0][19] ) );
  DFFASX1 \R_reg[0][18]  ( .D(n3190), .CLK(clk), .SETB(reset_n), .Q(\R[0][18] ) );
  DFFASX1 \R_reg[0][17]  ( .D(n3189), .CLK(clk), .SETB(reset_n), .Q(\R[0][17] ) );
  DFFASX1 \R_reg[0][16]  ( .D(n3188), .CLK(clk), .SETB(reset_n), .Q(\R[0][16] ) );
  DFFASX1 \R_reg[0][15]  ( .D(n3187), .CLK(clk), .SETB(reset_n), .Q(\R[0][15] ) );
  DFFASX1 \R_reg[0][14]  ( .D(n3186), .CLK(clk), .SETB(reset_n), .Q(\R[0][14] ) );
  DFFASX1 \R_reg[0][13]  ( .D(n3185), .CLK(clk), .SETB(reset_n), .Q(\R[0][13] ) );
  DFFASX1 \R_reg[0][12]  ( .D(n3184), .CLK(clk), .SETB(reset_n), .Q(\R[0][12] ) );
  DFFASX1 \R_reg[0][11]  ( .D(n3183), .CLK(clk), .SETB(reset_n), .Q(\R[0][11] ) );
  DFFASX1 \R_reg[0][10]  ( .D(n3182), .CLK(clk), .SETB(reset_n), .Q(\R[0][10] ) );
  DFFASX1 \R_reg[0][9]  ( .D(n3181), .CLK(clk), .SETB(reset_n), .Q(\R[0][9] )
         );
  DFFASX1 \R_reg[0][8]  ( .D(n3180), .CLK(clk), .SETB(reset_n), .Q(\R[0][8] )
         );
  DFFASX1 \R_reg[0][7]  ( .D(n3179), .CLK(clk), .SETB(reset_n), .Q(\R[0][7] )
         );
  DFFASX1 \R_reg[0][6]  ( .D(n3178), .CLK(clk), .SETB(reset_n), .Q(\R[0][6] )
         );
  DFFASX1 \R_reg[0][5]  ( .D(n3177), .CLK(clk), .SETB(reset_n), .Q(\R[0][5] )
         );
  DFFASX1 \R_reg[0][4]  ( .D(n3176), .CLK(clk), .SETB(reset_n), .Q(\R[0][4] )
         );
  DFFASX1 \R_reg[0][3]  ( .D(n3175), .CLK(clk), .SETB(reset_n), .Q(\R[0][3] )
         );
  DFFASX1 \R_reg[0][2]  ( .D(n3174), .CLK(clk), .SETB(reset_n), .Q(\R[0][2] )
         );
  DFFASX1 \R_reg[0][1]  ( .D(n3173), .CLK(clk), .SETB(reset_n), .Q(\R[0][1] )
         );
  DFFASX1 \R_reg[0][0]  ( .D(n3172), .CLK(clk), .SETB(reset_n), .Q(\R[0][0] )
         );
  thumb_DW01_addsub_0 r151 ( .A({1'b0, \U3/U74/Z_31 , \U3/U74/Z_30 , 
        \U3/U74/Z_29 , \U3/U74/Z_28 , \U3/U74/Z_27 , \U3/U74/Z_26 , 
        \U3/U74/Z_25 , \U3/U74/Z_24 , \U3/U74/Z_23 , \U3/U74/Z_22 , 
        \U3/U74/Z_21 , \U3/U74/Z_20 , \U3/U74/Z_19 , \U3/U74/Z_18 , 
        \U3/U74/Z_17 , \U3/U74/Z_16 , \U3/U74/Z_15 , \U3/U74/Z_14 , 
        \U3/U74/Z_13 , \U3/U74/Z_12 , \U3/U74/Z_11 , \U3/U74/Z_10 , 
        \U3/U74/Z_9 , \U3/U74/Z_8 , \U3/U74/Z_7 , \U3/U74/Z_6 , \U3/U74/Z_5 , 
        \U3/U74/Z_4 , \U3/U74/Z_3 , \U3/U74/Z_2 , \U3/U74/Z_1 , \U3/U74/Z_0 }), 
        .B({1'b0, \U3/U75/Z_31 , \U3/U75/Z_30 , \U3/U75/Z_29 , \U3/U75/Z_28 , 
        \U3/U75/Z_27 , \U3/U75/Z_26 , \U3/U75/Z_25 , \U3/U75/Z_24 , 
        \U3/U75/Z_23 , \U3/U75/Z_22 , \U3/U75/Z_21 , \U3/U75/Z_20 , 
        \U3/U75/Z_19 , \U3/U75/Z_18 , \U3/U75/Z_17 , \U3/U75/Z_16 , 
        \U3/U75/Z_15 , \U3/U75/Z_14 , \U3/U75/Z_13 , \U3/U75/Z_12 , 
        \U3/U75/Z_11 , \U3/U75/Z_10 , \U3/U75/Z_9 , \U3/U75/Z_8 , \U3/U75/Z_7 , 
        \U3/U75/Z_6 , \U3/U75/Z_5 , \U3/U75/Z_4 , \U3/U75/Z_3 , \U3/U75/Z_2 , 
        \U3/U75/Z_1 , \U3/U75/Z_0 }), .CI(\U3/U76/Z_0 ), .ADD_SUB(\U3/U77/Z_0 ), .SUM({n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
        n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
        n306, n307, n308, n309, n310, n311, n312, n313, n314}) );
  thumb_DW01_add_0 r1040 ( .A({1'b0, ID_Rn}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        ID_imm_offset[4:0], 1'b0, 1'b0}), .CI(1'b0), .SUM({N3588, N3587, N3586, 
        N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, 
        N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, 
        N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556})
         );
  thumb_DW01_add_1 r975 ( .A({1'b0, SP}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, ID_imm_offset, 1'b0, 1'b0}), .CI(
        1'b0), .SUM({N3687, N1244, N1243, N1242, N1241, N1240, N1239, N1238, 
        N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, 
        N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, 
        N1217, N1216, N1215, N1214, N1213}) );
  thumb_DW01_add_2 r974 ( .A({1'b0, ID_PC[31:2], 1'b0, 1'b0}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, ID_imm_offset, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N3654, N1212, N1211, N1210, N1209, 
        N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, 
        N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, 
        N1188, N1187, N1186, N1185, N1184, N1183, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}) );
  thumb_DW01_add_3 r973 ( .A({1'b0, ID_Rn}), .B({1'b0, N2429, ID_Rm_Rs[30:0]}), 
        .CI(1'b0), .SUM({N1180, N1179, N1178, N1177, N1176, N1175, N1174, 
        N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, 
        N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, 
        N1153, N1152, N1151, N1150, N1149, N1148}) );
  thumb_DW01_add_4 r969 ( .A(instruction_address), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0}), .CI(1'b0), .SUM({N232, N231, N230, N229, 
        N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, 
        N204, N203, N202, N201}) );
  thumb_DW_leftsh_2 sll_409 ( .A({1'b0, N2429, ID_Rm_Rs[30:0]}), .SH(
        ID_imm_offset[4:0]), .B({N3720, N3719, N3718, N3717, N3716, N3715, 
        N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, 
        N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, 
        N3694, N3693, N3692, N3691, N3690, N3689, N3688}) );
  thumb_DW_rightsh_2 srl_414 ( .A({N2429, ID_Rm_Rs[30:0], 1'b0}), .DATA_TC(
        1'b0), .SH(ID_imm_offset[4:0]), .B({N3822, N3821, N3820, N3819, N3818, 
        N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, 
        N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, 
        N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790}) );
  thumb_DW_rightsh_3 srl_417 ( .A({ID_Rd, 1'b0}), .DATA_TC(1'b0), .SH(
        ID_Rm_Rs[7:0]), .B({N3858, N3857, N3856, N3855, N3854, N3853, N3852, 
        N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, 
        N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, 
        N3831, N3830, N3829, N3828, N3827, N3826}) );
  thumb_DW_leftsh_3 sll_411 ( .A({1'b0, ID_Rd}), .SH(ID_Rm_Rs[7:0]), .B({N3756, 
        N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, 
        N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, 
        N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, 
        N3725, N3724}) );
  BSLEX1 \data_tri[0]  ( .INOUT1(n5740), .ENB(n5735), .INOUT2(data[0]) );
  BSLEX1 \data_tri[1]  ( .INOUT1(n5741), .ENB(n5735), .INOUT2(data[1]) );
  BSLEX1 \data_tri[2]  ( .INOUT1(n5742), .ENB(n5735), .INOUT2(data[2]) );
  BSLEX1 \data_tri[3]  ( .INOUT1(n5743), .ENB(n5735), .INOUT2(data[3]) );
  BSLEX1 \data_tri[4]  ( .INOUT1(n5744), .ENB(n5735), .INOUT2(data[4]) );
  BSLEX1 \data_tri[5]  ( .INOUT1(n5745), .ENB(n5735), .INOUT2(data[5]) );
  BSLEX1 \data_tri[6]  ( .INOUT1(n5746), .ENB(n5735), .INOUT2(data[6]) );
  BSLEX1 \data_tri[7]  ( .INOUT1(n5747), .ENB(n5735), .INOUT2(data[7]) );
  BSLEX1 \data_tri[8]  ( .INOUT1(n5748), .ENB(n5735), .INOUT2(data[8]) );
  BSLEX1 \data_tri[9]  ( .INOUT1(n5749), .ENB(n5735), .INOUT2(data[9]) );
  BSLEX1 \data_tri[10]  ( .INOUT1(n5750), .ENB(n5735), .INOUT2(data[10]) );
  BSLEX1 \data_tri[11]  ( .INOUT1(n5751), .ENB(n5735), .INOUT2(data[11]) );
  BSLEX1 \data_tri[12]  ( .INOUT1(n5752), .ENB(n5735), .INOUT2(data[12]) );
  BSLEX1 \data_tri[13]  ( .INOUT1(n5753), .ENB(n5735), .INOUT2(data[13]) );
  BSLEX1 \data_tri[14]  ( .INOUT1(n5754), .ENB(n5735), .INOUT2(data[14]) );
  BSLEX1 \data_tri[15]  ( .INOUT1(n5755), .ENB(n5735), .INOUT2(data[15]) );
  BSLEX1 \data_tri[16]  ( .INOUT1(n5756), .ENB(n5735), .INOUT2(data[16]) );
  BSLEX1 \data_tri[17]  ( .INOUT1(n5757), .ENB(n5735), .INOUT2(data[17]) );
  BSLEX1 \data_tri[18]  ( .INOUT1(n5758), .ENB(n5735), .INOUT2(data[18]) );
  BSLEX1 \data_tri[19]  ( .INOUT1(n5759), .ENB(n5735), .INOUT2(data[19]) );
  BSLEX1 \data_tri[20]  ( .INOUT1(n5760), .ENB(n5735), .INOUT2(data[20]) );
  BSLEX1 \data_tri[21]  ( .INOUT1(n5761), .ENB(n5735), .INOUT2(data[21]) );
  BSLEX1 \data_tri[22]  ( .INOUT1(n5762), .ENB(n5735), .INOUT2(data[22]) );
  BSLEX1 \data_tri[23]  ( .INOUT1(n5763), .ENB(n5735), .INOUT2(data[23]) );
  BSLEX1 \data_tri[24]  ( .INOUT1(n5764), .ENB(n5735), .INOUT2(data[24]) );
  BSLEX1 \data_tri[25]  ( .INOUT1(n5765), .ENB(n5735), .INOUT2(data[25]) );
  BSLEX1 \data_tri[26]  ( .INOUT1(n5766), .ENB(n5735), .INOUT2(data[26]) );
  BSLEX1 \data_tri[27]  ( .INOUT1(n5767), .ENB(n5735), .INOUT2(data[27]) );
  BSLEX1 \data_tri[28]  ( .INOUT1(n5768), .ENB(n5735), .INOUT2(data[28]) );
  BSLEX1 \data_tri[29]  ( .INOUT1(n5769), .ENB(n5735), .INOUT2(data[29]) );
  BSLEX1 \data_tri[30]  ( .INOUT1(n5770), .ENB(n5735), .INOUT2(data[30]) );
  BSLEX1 \data_tri[31]  ( .INOUT1(n5771), .ENB(n5735), .INOUT2(data[31]) );
  DFFX2 \ID_imm_offset_reg[1]  ( .D(n3632), .CLK(clk), .Q(ID_imm_offset[1]), 
        .QN(n2991) );
  DFFX2 \ID_imm_offset_reg[0]  ( .D(n3628), .CLK(clk), .Q(ID_imm_offset[0]), 
        .QN(n2988) );
  DFFX2 \ID_imm_offset_reg[2]  ( .D(n3636), .CLK(clk), .Q(ID_imm_offset[2]), 
        .QN(n2994) );
  DFFX2 \ID_imm_offset_reg[3]  ( .D(n3638), .CLK(clk), .Q(ID_imm_offset[3]), 
        .QN(n2995) );
  NOR2X1 U2887 ( .IN1(n4400), .IN2(n5019), .QN(n4438) );
  INVX2 U2888 ( .INP(n5163), .ZN(n4753) );
  NAND3X1 U2889 ( .IN1(n5723), .IN2(n5056), .IN3(n5720), .QN(\U3/U77/Z_0 ) );
  NOR2X1 U2890 ( .IN1(n4253), .IN2(N4634), .QN(n4326) );
  NOR2X1 U2891 ( .IN1(n5020), .IN2(n4400), .QN(n4439) );
  INVX0 U2892 ( .INP(n5728), .ZN(n4151) );
  INVX0 U2893 ( .INP(n5728), .ZN(n4152) );
  INVX0 U2894 ( .INP(n5728), .ZN(n4154) );
  INVX0 U2895 ( .INP(n5728), .ZN(n4153) );
  INVX0 U2896 ( .INP(n5728), .ZN(n4156) );
  INVX0 U2897 ( .INP(n5728), .ZN(n4155) );
  INVX0 U2898 ( .INP(n5728), .ZN(n4158) );
  INVX0 U2899 ( .INP(n5728), .ZN(n4157) );
  INVX0 U2900 ( .INP(n5728), .ZN(n4160) );
  INVX0 U2901 ( .INP(n5728), .ZN(n4159) );
  MUX41X1 U2902 ( .IN1(\R[5][30] ), .IN3(\R[7][30] ), .IN2(\R[4][30] ), .IN4(
        \R[6][30] ), .S0(N190), .S1(n5731), .Q(n4079) );
  MUX41X1 U2903 ( .IN1(\R[5][28] ), .IN3(\R[7][28] ), .IN2(\R[4][28] ), .IN4(
        \R[6][28] ), .S0(N190), .S1(n5731), .Q(n4075) );
  MUX41X1 U2904 ( .IN1(\R[5][26] ), .IN3(\R[7][26] ), .IN2(\R[4][26] ), .IN4(
        \R[6][26] ), .S0(N190), .S1(n5731), .Q(n4071) );
  MUX41X1 U2905 ( .IN1(\R[5][24] ), .IN3(\R[7][24] ), .IN2(\R[4][24] ), .IN4(
        \R[6][24] ), .S0(N190), .S1(n5731), .Q(n4067) );
  MUX41X1 U2906 ( .IN1(\R[5][21] ), .IN3(\R[7][21] ), .IN2(\R[4][21] ), .IN4(
        \R[6][21] ), .S0(N190), .S1(n5731), .Q(n4061) );
  INVX0 U2907 ( .INP(n3800), .ZN(n4225) );
  MUX41X1 U2908 ( .IN1(\R[7][19] ), .IN3(\R[5][19] ), .IN2(\R[6][19] ), .IN4(
        \R[4][19] ), .S0(n5730), .S1(n5731), .Q(n4057) );
  INVX0 U2909 ( .INP(n3800), .ZN(n4226) );
  INVX0 U2910 ( .INP(n3800), .ZN(n4227) );
  MUX41X1 U2911 ( .IN1(\R[7][17] ), .IN3(\R[5][17] ), .IN2(\R[6][17] ), .IN4(
        \R[4][17] ), .S0(n5730), .S1(n5731), .Q(n4053) );
  MUX41X1 U2912 ( .IN1(\R[7][15] ), .IN3(\R[5][15] ), .IN2(\R[6][15] ), .IN4(
        \R[4][15] ), .S0(n5730), .S1(n5731), .Q(n4049) );
  MUX41X1 U2913 ( .IN1(\R[7][12] ), .IN3(\R[5][12] ), .IN2(\R[6][12] ), .IN4(
        \R[4][12] ), .S0(n5730), .S1(n5731), .Q(n4043) );
  MUX41X1 U2914 ( .IN1(\R[7][10] ), .IN3(\R[5][10] ), .IN2(\R[6][10] ), .IN4(
        \R[4][10] ), .S0(n5730), .S1(n5731), .Q(n4039) );
  INVX0 U2915 ( .INP(n3800), .ZN(n4228) );
  INVX0 U2916 ( .INP(n3800), .ZN(n4229) );
  MUX41X1 U2917 ( .IN1(\R[7][8] ), .IN3(\R[5][8] ), .IN2(\R[6][8] ), .IN4(
        \R[4][8] ), .S0(n5730), .S1(n5731), .Q(n4035) );
  INVX0 U2918 ( .INP(n3800), .ZN(n4230) );
  INVX0 U2919 ( .INP(n3800), .ZN(n4231) );
  MUX41X1 U2920 ( .IN1(\R[7][6] ), .IN3(\R[5][6] ), .IN2(\R[6][6] ), .IN4(
        \R[4][6] ), .S0(n5730), .S1(n5731), .Q(n4031) );
  INVX0 U2921 ( .INP(n3800), .ZN(n4232) );
  INVX0 U2922 ( .INP(n3800), .ZN(n4233) );
  MUX41X1 U2923 ( .IN1(\R[7][4] ), .IN3(\R[5][4] ), .IN2(\R[6][4] ), .IN4(
        \R[4][4] ), .S0(n5730), .S1(n5731), .Q(n4027) );
  INVX0 U2924 ( .INP(n3800), .ZN(n4234) );
  INVX0 U2925 ( .INP(n3800), .ZN(n4235) );
  INVX0 U2926 ( .INP(n3800), .ZN(n4236) );
  MUX41X1 U2927 ( .IN1(\R[7][1] ), .IN3(\R[5][1] ), .IN2(\R[6][1] ), .IN4(
        \R[4][1] ), .S0(n5730), .S1(n5731), .Q(n4021) );
  INVX0 U2928 ( .INP(n3800), .ZN(n4237) );
  INVX0 U2929 ( .INP(n3800), .ZN(n4238) );
  MUX41X1 U2930 ( .IN1(\R[3][31] ), .IN3(\R[1][31] ), .IN2(\R[2][31] ), .IN4(
        \R[0][31] ), .S0(n5730), .S1(n5731), .Q(n4082) );
  MUX41X1 U2931 ( .IN1(\R[3][29] ), .IN3(\R[1][29] ), .IN2(\R[2][29] ), .IN4(
        \R[0][29] ), .S0(n5730), .S1(n5731), .Q(n4078) );
  MUX41X1 U2932 ( .IN1(\R[3][27] ), .IN3(\R[1][27] ), .IN2(\R[2][27] ), .IN4(
        \R[0][27] ), .S0(n5730), .S1(n5731), .Q(n4074) );
  MUX41X1 U2933 ( .IN1(\R[3][24] ), .IN3(\R[1][24] ), .IN2(\R[2][24] ), .IN4(
        \R[0][24] ), .S0(n5730), .S1(n5731), .Q(n4068) );
  MUX41X1 U2934 ( .IN1(\R[3][22] ), .IN3(\R[1][22] ), .IN2(\R[2][22] ), .IN4(
        \R[0][22] ), .S0(n5730), .S1(n5731), .Q(n4064) );
  MUX41X1 U2935 ( .IN1(\R[3][20] ), .IN3(\R[1][20] ), .IN2(\R[2][20] ), .IN4(
        \R[0][20] ), .S0(n5730), .S1(n5731), .Q(n4060) );
  MUX41X1 U2936 ( .IN1(\R[3][18] ), .IN3(\R[1][18] ), .IN2(\R[2][18] ), .IN4(
        \R[0][18] ), .S0(n5730), .S1(n5731), .Q(n4056) );
  MUX41X1 U2937 ( .IN1(\R[3][16] ), .IN3(\R[1][16] ), .IN2(\R[2][16] ), .IN4(
        \R[0][16] ), .S0(n5730), .S1(n5731), .Q(n4052) );
  MUX41X1 U2938 ( .IN1(\R[3][13] ), .IN3(\R[1][13] ), .IN2(\R[2][13] ), .IN4(
        \R[0][13] ), .S0(n5730), .S1(n5731), .Q(n4046) );
  INVX0 U2939 ( .INP(n5731), .ZN(n4083) );
  INVX0 U2940 ( .INP(n5731), .ZN(n4084) );
  INVX0 U2941 ( .INP(n5731), .ZN(n4085) );
  INVX0 U2942 ( .INP(n5731), .ZN(n4086) );
  MUX41X1 U2943 ( .IN1(\R[3][31] ), .IN3(\R[1][31] ), .IN2(\R[2][31] ), .IN4(
        \R[0][31] ), .S0(n5733), .S1(n5734), .Q(n4011) );
  MUX41X1 U2944 ( .IN1(\R[3][29] ), .IN3(\R[1][29] ), .IN2(\R[2][29] ), .IN4(
        \R[0][29] ), .S0(n5733), .S1(n5734), .Q(n4007) );
  MUX41X1 U2945 ( .IN1(\R[3][27] ), .IN3(\R[1][27] ), .IN2(\R[2][27] ), .IN4(
        \R[0][27] ), .S0(n5733), .S1(n5734), .Q(n4003) );
  MUX41X1 U2946 ( .IN1(\R[3][24] ), .IN3(\R[1][24] ), .IN2(\R[2][24] ), .IN4(
        \R[0][24] ), .S0(n5733), .S1(n5734), .Q(n3997) );
  MUX41X1 U2947 ( .IN1(\R[3][22] ), .IN3(\R[1][22] ), .IN2(\R[2][22] ), .IN4(
        \R[0][22] ), .S0(n5733), .S1(n5734), .Q(n3993) );
  MUX41X1 U2948 ( .IN1(\R[3][20] ), .IN3(\R[1][20] ), .IN2(\R[2][20] ), .IN4(
        \R[0][20] ), .S0(n5733), .S1(n5734), .Q(n3989) );
  MUX41X1 U2949 ( .IN1(\R[3][18] ), .IN3(\R[1][18] ), .IN2(\R[2][18] ), .IN4(
        \R[0][18] ), .S0(n5733), .S1(n5734), .Q(n3985) );
  MUX41X1 U2950 ( .IN1(\R[3][16] ), .IN3(\R[1][16] ), .IN2(\R[2][16] ), .IN4(
        \R[0][16] ), .S0(n5733), .S1(n5734), .Q(n3981) );
  MUX41X1 U2951 ( .IN1(\R[3][13] ), .IN3(\R[1][13] ), .IN2(\R[2][13] ), .IN4(
        \R[0][13] ), .S0(n5733), .S1(n5734), .Q(n3975) );
  INVX0 U2952 ( .INP(n5734), .ZN(n4012) );
  INVX0 U2953 ( .INP(n5734), .ZN(n4013) );
  INVX0 U2954 ( .INP(n5734), .ZN(n4014) );
  INVX0 U2955 ( .INP(n5734), .ZN(n4015) );
  INVX0 U2956 ( .INP(n5734), .ZN(n4016) );
  INVX0 U2957 ( .INP(n5734), .ZN(n4017) );
  INVX0 U2958 ( .INP(n5734), .ZN(n4018) );
  XOR2X1 U2959 ( .IN1(n3132), .IN2(IF_IR[13]), .Q(n3918) );
  MUX21X1 U2960 ( .IN1(IF_IR[12]), .IN2(N690), .S(IF_IR[13]), .Q(n3919) );
  AND2X1 U2961 ( .IN1(N695), .IN2(n3130), .Q(n3920) );
  MUX21X1 U2962 ( .IN1(n3919), .IN2(n3920), .S(IF_IR[14]), .Q(n3921) );
  OR2X1 U2963 ( .IN1(n3795), .IN2(IF_IR[13]), .Q(n3922) );
  MUX21X1 U2964 ( .IN1(n3922), .IN2(n3947), .S(IF_IR[14]), .Q(n3923) );
  MUX21X1 U2965 ( .IN1(n3923), .IN2(n3921), .S(IF_IR[15]), .Q(N773) );
  OR2X1 U2966 ( .IN1(n5738), .IN2(IF_IR[13]), .Q(n3924) );
  MUX21X1 U2967 ( .IN1(n3924), .IN2(n3947), .S(IF_IR[14]), .Q(n3925) );
  MUX21X1 U2968 ( .IN1(n3925), .IN2(n3921), .S(IF_IR[15]), .Q(N777) );
  MUX21X1 U2969 ( .IN1(n3799), .IN2(N693), .S(IF_IR[14]), .Q(n3926) );
  OR2X1 U2970 ( .IN1(N688), .IN2(IF_IR[14]), .Q(n3927) );
  MUX21X1 U2971 ( .IN1(n5737), .IN2(n3799), .S(IF_IR[14]), .Q(n3928) );
  MUX21X1 U2972 ( .IN1(N550), .IN2(N599), .S(IF_IR[14]), .Q(n3929) );
  MUX41X1 U2973 ( .IN1(n3929), .IN3(n3928), .IN2(n3926), .IN4(n3927), .S0(
        IF_IR[13]), .S1(IF_IR[15]), .Q(N772) );
  MUX21X1 U2974 ( .IN1(N693), .IN2(N688), .S(IF_IR[13]), .Q(n3930) );
  MUX21X1 U2975 ( .IN1(N548), .IN2(N598), .S(IF_IR[14]), .Q(n3931) );
  MUX21X1 U2976 ( .IN1(n3931), .IN2(IF_IR[11]), .S(IF_IR[13]), .Q(n3932) );
  OR2X1 U2977 ( .IN1(n3918), .IN2(n3930), .Q(n3933) );
  MUX21X1 U2978 ( .IN1(n3932), .IN2(n3933), .S(IF_IR[15]), .Q(N771) );
  MUX21X1 U2979 ( .IN1(IF_IR[11]), .IN2(N687), .S(IF_IR[15]), .Q(n3934) );
  MUX41X1 U2980 ( .IN1(N548), .IN3(N596), .IN2(IF_IR[11]), .IN4(n5736), .S0(
        IF_IR[14]), .S1(IF_IR[15]), .Q(n3935) );
  OR2X1 U2981 ( .IN1(IF_IR[14]), .IN2(n3934), .Q(n3936) );
  MUX21X1 U2982 ( .IN1(n3935), .IN2(n3936), .S(IF_IR[13]), .Q(N769) );
  MUX21X1 U2983 ( .IN1(IF_IR[11]), .IN2(N694), .S(IF_IR[14]), .Q(n3937) );
  OR2X1 U2984 ( .IN1(N686), .IN2(IF_IR[14]), .Q(n3938) );
  MUX21X1 U2985 ( .IN1(N547), .IN2(N595), .S(IF_IR[14]), .Q(n3939) );
  OR2X1 U2986 ( .IN1(n3799), .IN2(n3132), .Q(n3940) );
  MUX41X1 U2987 ( .IN1(n3939), .IN3(n3940), .IN2(n3937), .IN4(n3938), .S0(
        IF_IR[13]), .S1(IF_IR[15]), .Q(N768) );
  MUX21X1 U2988 ( .IN1(IF_IR[11]), .IN2(N693), .S(IF_IR[14]), .Q(n3941) );
  OR2X1 U2989 ( .IN1(N685), .IN2(IF_IR[14]), .Q(n3942) );
  MUX21X1 U2990 ( .IN1(n3941), .IN2(n3942), .S(IF_IR[13]), .Q(n3943) );
  AND2X1 U2991 ( .IN1(n3945), .IN2(n3130), .Q(n3944) );
  MUX21X1 U2992 ( .IN1(n3944), .IN2(n3943), .S(IF_IR[15]), .Q(N767) );
  MUX21X1 U2993 ( .IN1(n5739), .IN2(IF_IR[12]), .S(IF_IR[13]), .Q(n3946) );
  MUX21X1 U2994 ( .IN1(N498), .IN2(n5739), .S(IF_IR[14]), .Q(n3945) );
  INVX0 U2995 ( .INP(n3946), .ZN(n3947) );
  MUX41X1 U2996 ( .IN1(\R[4][0] ), .IN3(\R[6][0] ), .IN2(\R[5][0] ), .IN4(
        \R[7][0] ), .S0(N187), .S1(n4012), .Q(n3948) );
  MUX41X1 U2997 ( .IN1(\R[0][0] ), .IN3(\R[2][0] ), .IN2(\R[1][0] ), .IN4(
        \R[3][0] ), .S0(N187), .S1(n4012), .Q(n3949) );
  MUX21X1 U2998 ( .IN1(n3949), .IN2(n3948), .S(N188), .Q(N376) );
  MUX41X1 U2999 ( .IN1(\R[4][1] ), .IN3(\R[6][1] ), .IN2(\R[5][1] ), .IN4(
        \R[7][1] ), .S0(N187), .S1(n4015), .Q(n3950) );
  MUX41X1 U3000 ( .IN1(\R[0][1] ), .IN3(\R[2][1] ), .IN2(\R[1][1] ), .IN4(
        \R[3][1] ), .S0(N187), .S1(n4017), .Q(n3951) );
  MUX21X1 U3001 ( .IN1(n3951), .IN2(n3950), .S(N188), .Q(N375) );
  MUX41X1 U3002 ( .IN1(\R[4][2] ), .IN3(\R[6][2] ), .IN2(\R[5][2] ), .IN4(
        \R[7][2] ), .S0(N187), .S1(n4015), .Q(n3952) );
  MUX41X1 U3003 ( .IN1(\R[0][2] ), .IN3(\R[2][2] ), .IN2(\R[1][2] ), .IN4(
        \R[3][2] ), .S0(N187), .S1(n4018), .Q(n3953) );
  MUX21X1 U3004 ( .IN1(n3953), .IN2(n3952), .S(N188), .Q(N374) );
  MUX41X1 U3005 ( .IN1(\R[4][3] ), .IN3(\R[6][3] ), .IN2(\R[5][3] ), .IN4(
        \R[7][3] ), .S0(N187), .S1(n4016), .Q(n3954) );
  MUX41X1 U3006 ( .IN1(\R[0][3] ), .IN3(\R[2][3] ), .IN2(\R[1][3] ), .IN4(
        \R[3][3] ), .S0(N187), .S1(n4017), .Q(n3955) );
  MUX21X1 U3007 ( .IN1(n3955), .IN2(n3954), .S(N188), .Q(N373) );
  MUX41X1 U3008 ( .IN1(\R[4][4] ), .IN3(\R[6][4] ), .IN2(\R[5][4] ), .IN4(
        \R[7][4] ), .S0(N187), .S1(n4013), .Q(n3956) );
  MUX41X1 U3009 ( .IN1(\R[0][4] ), .IN3(\R[2][4] ), .IN2(\R[1][4] ), .IN4(
        \R[3][4] ), .S0(N187), .S1(n4016), .Q(n3957) );
  MUX21X1 U3010 ( .IN1(n3957), .IN2(n3956), .S(N188), .Q(N372) );
  MUX41X1 U3011 ( .IN1(\R[4][5] ), .IN3(\R[6][5] ), .IN2(\R[5][5] ), .IN4(
        \R[7][5] ), .S0(N187), .S1(n4018), .Q(n3958) );
  MUX41X1 U3012 ( .IN1(\R[0][5] ), .IN3(\R[2][5] ), .IN2(\R[1][5] ), .IN4(
        \R[3][5] ), .S0(N187), .S1(n4015), .Q(n3959) );
  MUX21X1 U3013 ( .IN1(n3959), .IN2(n3958), .S(N188), .Q(N371) );
  MUX41X1 U3014 ( .IN1(\R[4][6] ), .IN3(\R[6][6] ), .IN2(\R[5][6] ), .IN4(
        \R[7][6] ), .S0(N187), .S1(n4012), .Q(n3960) );
  MUX41X1 U3015 ( .IN1(\R[0][6] ), .IN3(\R[2][6] ), .IN2(\R[1][6] ), .IN4(
        \R[3][6] ), .S0(N187), .S1(n4014), .Q(n3961) );
  MUX21X1 U3016 ( .IN1(n3961), .IN2(n3960), .S(N188), .Q(N370) );
  MUX41X1 U3017 ( .IN1(\R[4][7] ), .IN3(\R[6][7] ), .IN2(\R[5][7] ), .IN4(
        \R[7][7] ), .S0(N187), .S1(n4018), .Q(n3962) );
  MUX41X1 U3018 ( .IN1(\R[0][7] ), .IN3(\R[2][7] ), .IN2(\R[1][7] ), .IN4(
        \R[3][7] ), .S0(N187), .S1(n4013), .Q(n3963) );
  MUX21X1 U3019 ( .IN1(n3963), .IN2(n3962), .S(N188), .Q(N369) );
  MUX41X1 U3020 ( .IN1(\R[4][8] ), .IN3(\R[6][8] ), .IN2(\R[5][8] ), .IN4(
        \R[7][8] ), .S0(N187), .S1(n5718), .Q(n3964) );
  MUX41X1 U3021 ( .IN1(\R[0][8] ), .IN3(\R[2][8] ), .IN2(\R[1][8] ), .IN4(
        \R[3][8] ), .S0(N187), .S1(n4012), .Q(n3965) );
  MUX21X1 U3022 ( .IN1(n3965), .IN2(n3964), .S(N188), .Q(N368) );
  MUX41X1 U3023 ( .IN1(\R[4][9] ), .IN3(\R[6][9] ), .IN2(\R[5][9] ), .IN4(
        \R[7][9] ), .S0(N187), .S1(n4016), .Q(n3966) );
  MUX41X1 U3024 ( .IN1(\R[0][9] ), .IN3(\R[2][9] ), .IN2(\R[1][9] ), .IN4(
        \R[3][9] ), .S0(N187), .S1(n4018), .Q(n3967) );
  MUX21X1 U3025 ( .IN1(n3967), .IN2(n3966), .S(N188), .Q(N367) );
  MUX41X1 U3026 ( .IN1(\R[4][10] ), .IN3(\R[6][10] ), .IN2(\R[5][10] ), .IN4(
        \R[7][10] ), .S0(N187), .S1(n4018), .Q(n3968) );
  MUX41X1 U3027 ( .IN1(\R[0][10] ), .IN3(\R[2][10] ), .IN2(\R[1][10] ), .IN4(
        \R[3][10] ), .S0(N187), .S1(n4015), .Q(n3969) );
  MUX21X1 U3028 ( .IN1(n3969), .IN2(n3968), .S(N188), .Q(N366) );
  MUX41X1 U3029 ( .IN1(\R[4][11] ), .IN3(\R[6][11] ), .IN2(\R[5][11] ), .IN4(
        \R[7][11] ), .S0(N187), .S1(n4014), .Q(n3970) );
  MUX41X1 U3030 ( .IN1(\R[0][11] ), .IN3(\R[2][11] ), .IN2(\R[1][11] ), .IN4(
        \R[3][11] ), .S0(N187), .S1(n4013), .Q(n3971) );
  MUX21X1 U3031 ( .IN1(n3971), .IN2(n3970), .S(N188), .Q(N365) );
  MUX41X1 U3032 ( .IN1(\R[4][12] ), .IN3(\R[6][12] ), .IN2(\R[5][12] ), .IN4(
        \R[7][12] ), .S0(N187), .S1(n4015), .Q(n3972) );
  MUX41X1 U3033 ( .IN1(\R[0][12] ), .IN3(\R[2][12] ), .IN2(\R[1][12] ), .IN4(
        \R[3][12] ), .S0(N187), .S1(n4014), .Q(n3973) );
  MUX21X1 U3034 ( .IN1(n3973), .IN2(n3972), .S(N188), .Q(N364) );
  MUX41X1 U3035 ( .IN1(\R[4][13] ), .IN3(\R[6][13] ), .IN2(\R[5][13] ), .IN4(
        \R[7][13] ), .S0(N187), .S1(n4017), .Q(n3974) );
  MUX21X1 U3036 ( .IN1(n3975), .IN2(n3974), .S(N188), .Q(N363) );
  MUX41X1 U3037 ( .IN1(\R[4][14] ), .IN3(\R[6][14] ), .IN2(\R[5][14] ), .IN4(
        \R[7][14] ), .S0(N187), .S1(n5718), .Q(n3976) );
  MUX41X1 U3038 ( .IN1(\R[0][14] ), .IN3(\R[2][14] ), .IN2(\R[1][14] ), .IN4(
        \R[3][14] ), .S0(N187), .S1(n5718), .Q(n3977) );
  MUX21X1 U3039 ( .IN1(n3977), .IN2(n3976), .S(N188), .Q(N362) );
  MUX41X1 U3040 ( .IN1(\R[4][15] ), .IN3(\R[6][15] ), .IN2(\R[5][15] ), .IN4(
        \R[7][15] ), .S0(N187), .S1(n4012), .Q(n3978) );
  MUX41X1 U3041 ( .IN1(\R[0][15] ), .IN3(\R[2][15] ), .IN2(\R[1][15] ), .IN4(
        \R[3][15] ), .S0(N187), .S1(n4017), .Q(n3979) );
  MUX21X1 U3042 ( .IN1(n3979), .IN2(n3978), .S(N188), .Q(N361) );
  MUX41X1 U3043 ( .IN1(\R[4][16] ), .IN3(\R[6][16] ), .IN2(\R[5][16] ), .IN4(
        \R[7][16] ), .S0(N187), .S1(n4017), .Q(n3980) );
  MUX21X1 U3044 ( .IN1(n3981), .IN2(n3980), .S(N188), .Q(N360) );
  MUX41X1 U3045 ( .IN1(\R[4][17] ), .IN3(\R[6][17] ), .IN2(\R[5][17] ), .IN4(
        \R[7][17] ), .S0(N187), .S1(n4015), .Q(n3982) );
  MUX41X1 U3046 ( .IN1(\R[0][17] ), .IN3(\R[2][17] ), .IN2(\R[1][17] ), .IN4(
        \R[3][17] ), .S0(N187), .S1(n4014), .Q(n3983) );
  MUX21X1 U3047 ( .IN1(n3983), .IN2(n3982), .S(N188), .Q(N359) );
  MUX41X1 U3048 ( .IN1(\R[4][18] ), .IN3(\R[6][18] ), .IN2(\R[5][18] ), .IN4(
        \R[7][18] ), .S0(N187), .S1(n4013), .Q(n3984) );
  MUX21X1 U3049 ( .IN1(n3985), .IN2(n3984), .S(N188), .Q(N358) );
  MUX41X1 U3050 ( .IN1(\R[4][19] ), .IN3(\R[6][19] ), .IN2(\R[5][19] ), .IN4(
        \R[7][19] ), .S0(N187), .S1(n4016), .Q(n3986) );
  MUX41X1 U3051 ( .IN1(\R[0][19] ), .IN3(\R[2][19] ), .IN2(\R[1][19] ), .IN4(
        \R[3][19] ), .S0(N187), .S1(n4013), .Q(n3987) );
  MUX21X1 U3052 ( .IN1(n3987), .IN2(n3986), .S(N188), .Q(N357) );
  MUX41X1 U3053 ( .IN1(\R[4][20] ), .IN3(\R[6][20] ), .IN2(\R[5][20] ), .IN4(
        \R[7][20] ), .S0(N187), .S1(n5718), .Q(n3988) );
  MUX21X1 U3054 ( .IN1(n3989), .IN2(n3988), .S(N188), .Q(N356) );
  MUX41X1 U3055 ( .IN1(\R[4][21] ), .IN3(\R[6][21] ), .IN2(\R[5][21] ), .IN4(
        \R[7][21] ), .S0(N187), .S1(n4013), .Q(n3990) );
  MUX41X1 U3056 ( .IN1(\R[0][21] ), .IN3(\R[2][21] ), .IN2(\R[1][21] ), .IN4(
        \R[3][21] ), .S0(N187), .S1(n4017), .Q(n3991) );
  MUX21X1 U3057 ( .IN1(n3991), .IN2(n3990), .S(N188), .Q(N355) );
  MUX41X1 U3058 ( .IN1(\R[4][22] ), .IN3(\R[6][22] ), .IN2(\R[5][22] ), .IN4(
        \R[7][22] ), .S0(N187), .S1(n4012), .Q(n3992) );
  MUX21X1 U3059 ( .IN1(n3993), .IN2(n3992), .S(N188), .Q(N354) );
  MUX41X1 U3060 ( .IN1(\R[4][23] ), .IN3(\R[6][23] ), .IN2(\R[5][23] ), .IN4(
        \R[7][23] ), .S0(N187), .S1(n4018), .Q(n3994) );
  MUX41X1 U3061 ( .IN1(\R[0][23] ), .IN3(\R[2][23] ), .IN2(\R[1][23] ), .IN4(
        \R[3][23] ), .S0(N187), .S1(n4017), .Q(n3995) );
  MUX21X1 U3062 ( .IN1(n3995), .IN2(n3994), .S(N188), .Q(N353) );
  MUX41X1 U3063 ( .IN1(\R[4][24] ), .IN3(\R[6][24] ), .IN2(\R[5][24] ), .IN4(
        \R[7][24] ), .S0(N187), .S1(n4016), .Q(n3996) );
  MUX21X1 U3064 ( .IN1(n3997), .IN2(n3996), .S(N188), .Q(N352) );
  MUX41X1 U3065 ( .IN1(\R[4][25] ), .IN3(\R[6][25] ), .IN2(\R[5][25] ), .IN4(
        \R[7][25] ), .S0(N187), .S1(n4016), .Q(n3998) );
  MUX41X1 U3066 ( .IN1(\R[0][25] ), .IN3(\R[2][25] ), .IN2(\R[1][25] ), .IN4(
        \R[3][25] ), .S0(N187), .S1(n4014), .Q(n3999) );
  MUX21X1 U3067 ( .IN1(n3999), .IN2(n3998), .S(N188), .Q(N351) );
  MUX41X1 U3068 ( .IN1(\R[4][26] ), .IN3(\R[6][26] ), .IN2(\R[5][26] ), .IN4(
        \R[7][26] ), .S0(N187), .S1(n5718), .Q(n4000) );
  MUX41X1 U3069 ( .IN1(\R[0][26] ), .IN3(\R[2][26] ), .IN2(\R[1][26] ), .IN4(
        \R[3][26] ), .S0(N187), .S1(n4014), .Q(n4001) );
  MUX21X1 U3070 ( .IN1(n4001), .IN2(n4000), .S(N188), .Q(N350) );
  MUX41X1 U3071 ( .IN1(\R[4][27] ), .IN3(\R[6][27] ), .IN2(\R[5][27] ), .IN4(
        \R[7][27] ), .S0(N187), .S1(n4012), .Q(n4002) );
  MUX21X1 U3072 ( .IN1(n4003), .IN2(n4002), .S(N188), .Q(N349) );
  MUX41X1 U3073 ( .IN1(\R[4][28] ), .IN3(\R[6][28] ), .IN2(\R[5][28] ), .IN4(
        \R[7][28] ), .S0(N187), .S1(n4014), .Q(n4004) );
  MUX41X1 U3074 ( .IN1(\R[0][28] ), .IN3(\R[2][28] ), .IN2(\R[1][28] ), .IN4(
        \R[3][28] ), .S0(N187), .S1(n4018), .Q(n4005) );
  MUX21X1 U3075 ( .IN1(n4005), .IN2(n4004), .S(N188), .Q(N348) );
  MUX41X1 U3076 ( .IN1(\R[4][29] ), .IN3(\R[6][29] ), .IN2(\R[5][29] ), .IN4(
        \R[7][29] ), .S0(N187), .S1(n4013), .Q(n4006) );
  MUX21X1 U3077 ( .IN1(n4007), .IN2(n4006), .S(N188), .Q(N347) );
  MUX41X1 U3078 ( .IN1(\R[4][30] ), .IN3(\R[6][30] ), .IN2(\R[5][30] ), .IN4(
        \R[7][30] ), .S0(N187), .S1(n4016), .Q(n4008) );
  MUX41X1 U3079 ( .IN1(\R[0][30] ), .IN3(\R[2][30] ), .IN2(\R[1][30] ), .IN4(
        \R[3][30] ), .S0(N187), .S1(n4015), .Q(n4009) );
  MUX21X1 U3080 ( .IN1(n4009), .IN2(n4008), .S(N188), .Q(N346) );
  MUX41X1 U3081 ( .IN1(\R[4][31] ), .IN3(\R[6][31] ), .IN2(\R[5][31] ), .IN4(
        \R[7][31] ), .S0(N187), .S1(n5718), .Q(n4010) );
  MUX21X1 U3082 ( .IN1(n4011), .IN2(n4010), .S(N188), .Q(N345) );
  MUX41X1 U3083 ( .IN1(\R[4][0] ), .IN3(\R[6][0] ), .IN2(\R[5][0] ), .IN4(
        \R[7][0] ), .S0(N190), .S1(n4086), .Q(n4019) );
  MUX41X1 U3084 ( .IN1(\R[0][0] ), .IN3(\R[2][0] ), .IN2(\R[1][0] ), .IN4(
        \R[3][0] ), .S0(N190), .S1(n4084), .Q(n4020) );
  MUX21X1 U3085 ( .IN1(n4020), .IN2(n4019), .S(N191), .Q(N408) );
  MUX41X1 U3086 ( .IN1(\R[0][1] ), .IN3(\R[2][1] ), .IN2(\R[1][1] ), .IN4(
        \R[3][1] ), .S0(N190), .S1(n4086), .Q(n4022) );
  MUX21X1 U3087 ( .IN1(n4022), .IN2(n4021), .S(N191), .Q(N407) );
  MUX41X1 U3088 ( .IN1(\R[4][2] ), .IN3(\R[6][2] ), .IN2(\R[5][2] ), .IN4(
        \R[7][2] ), .S0(N190), .S1(n4085), .Q(n4023) );
  MUX41X1 U3089 ( .IN1(\R[0][2] ), .IN3(\R[2][2] ), .IN2(\R[1][2] ), .IN4(
        \R[3][2] ), .S0(N190), .S1(n4085), .Q(n4024) );
  MUX21X1 U3090 ( .IN1(n4024), .IN2(n4023), .S(N191), .Q(N406) );
  MUX41X1 U3091 ( .IN1(\R[4][3] ), .IN3(\R[6][3] ), .IN2(\R[5][3] ), .IN4(
        \R[7][3] ), .S0(N190), .S1(n4086), .Q(n4025) );
  MUX41X1 U3092 ( .IN1(\R[0][3] ), .IN3(\R[2][3] ), .IN2(\R[1][3] ), .IN4(
        \R[3][3] ), .S0(N190), .S1(n4084), .Q(n4026) );
  MUX21X1 U3093 ( .IN1(n4026), .IN2(n4025), .S(N191), .Q(N405) );
  MUX41X1 U3094 ( .IN1(\R[0][4] ), .IN3(\R[2][4] ), .IN2(\R[1][4] ), .IN4(
        \R[3][4] ), .S0(N190), .S1(n4083), .Q(n4028) );
  MUX21X1 U3095 ( .IN1(n4028), .IN2(n4027), .S(N191), .Q(N404) );
  MUX41X1 U3096 ( .IN1(\R[4][5] ), .IN3(\R[6][5] ), .IN2(\R[5][5] ), .IN4(
        \R[7][5] ), .S0(N190), .S1(n4083), .Q(n4029) );
  MUX41X1 U3097 ( .IN1(\R[0][5] ), .IN3(\R[2][5] ), .IN2(\R[1][5] ), .IN4(
        \R[3][5] ), .S0(N190), .S1(n4085), .Q(n4030) );
  MUX21X1 U3098 ( .IN1(n4030), .IN2(n4029), .S(N191), .Q(N403) );
  MUX41X1 U3099 ( .IN1(\R[0][6] ), .IN3(\R[2][6] ), .IN2(\R[1][6] ), .IN4(
        \R[3][6] ), .S0(N190), .S1(n5715), .Q(n4032) );
  MUX21X1 U3100 ( .IN1(n4032), .IN2(n4031), .S(N191), .Q(N402) );
  MUX41X1 U3101 ( .IN1(\R[4][7] ), .IN3(\R[6][7] ), .IN2(\R[5][7] ), .IN4(
        \R[7][7] ), .S0(N190), .S1(n5715), .Q(n4033) );
  MUX41X1 U3102 ( .IN1(\R[0][7] ), .IN3(\R[2][7] ), .IN2(\R[1][7] ), .IN4(
        \R[3][7] ), .S0(N190), .S1(n4084), .Q(n4034) );
  MUX21X1 U3103 ( .IN1(n4034), .IN2(n4033), .S(N191), .Q(N401) );
  MUX41X1 U3104 ( .IN1(\R[0][8] ), .IN3(\R[2][8] ), .IN2(\R[1][8] ), .IN4(
        \R[3][8] ), .S0(N190), .S1(n4084), .Q(n4036) );
  MUX21X1 U3105 ( .IN1(n4036), .IN2(n4035), .S(N191), .Q(N400) );
  MUX41X1 U3106 ( .IN1(\R[4][9] ), .IN3(\R[6][9] ), .IN2(\R[5][9] ), .IN4(
        \R[7][9] ), .S0(N190), .S1(n4085), .Q(n4037) );
  MUX41X1 U3107 ( .IN1(\R[0][9] ), .IN3(\R[2][9] ), .IN2(\R[1][9] ), .IN4(
        \R[3][9] ), .S0(N190), .S1(n5715), .Q(n4038) );
  MUX21X1 U3108 ( .IN1(n4038), .IN2(n4037), .S(N191), .Q(N399) );
  MUX41X1 U3109 ( .IN1(\R[0][10] ), .IN3(\R[2][10] ), .IN2(\R[1][10] ), .IN4(
        \R[3][10] ), .S0(N190), .S1(n4086), .Q(n4040) );
  MUX21X1 U3110 ( .IN1(n4040), .IN2(n4039), .S(N191), .Q(N398) );
  MUX41X1 U3111 ( .IN1(\R[4][11] ), .IN3(\R[6][11] ), .IN2(\R[5][11] ), .IN4(
        \R[7][11] ), .S0(N190), .S1(n4084), .Q(n4041) );
  MUX41X1 U3112 ( .IN1(\R[0][11] ), .IN3(\R[2][11] ), .IN2(\R[1][11] ), .IN4(
        \R[3][11] ), .S0(N190), .S1(n4085), .Q(n4042) );
  MUX21X1 U3113 ( .IN1(n4042), .IN2(n4041), .S(N191), .Q(N397) );
  MUX41X1 U3114 ( .IN1(\R[0][12] ), .IN3(\R[2][12] ), .IN2(\R[1][12] ), .IN4(
        \R[3][12] ), .S0(N190), .S1(n4085), .Q(n4044) );
  MUX21X1 U3115 ( .IN1(n4044), .IN2(n4043), .S(N191), .Q(N396) );
  MUX41X1 U3116 ( .IN1(\R[4][13] ), .IN3(\R[6][13] ), .IN2(\R[5][13] ), .IN4(
        \R[7][13] ), .S0(N190), .S1(n5715), .Q(n4045) );
  MUX21X1 U3117 ( .IN1(n4046), .IN2(n4045), .S(N191), .Q(N395) );
  MUX41X1 U3118 ( .IN1(\R[4][14] ), .IN3(\R[6][14] ), .IN2(\R[5][14] ), .IN4(
        \R[7][14] ), .S0(N190), .S1(n4084), .Q(n4047) );
  MUX41X1 U3119 ( .IN1(\R[0][14] ), .IN3(\R[2][14] ), .IN2(\R[1][14] ), .IN4(
        \R[3][14] ), .S0(N190), .S1(n4083), .Q(n4048) );
  MUX21X1 U3120 ( .IN1(n4048), .IN2(n4047), .S(N191), .Q(N394) );
  MUX41X1 U3121 ( .IN1(\R[0][15] ), .IN3(\R[2][15] ), .IN2(\R[1][15] ), .IN4(
        \R[3][15] ), .S0(N190), .S1(n4086), .Q(n4050) );
  MUX21X1 U3122 ( .IN1(n4050), .IN2(n4049), .S(N191), .Q(N393) );
  MUX41X1 U3123 ( .IN1(\R[4][16] ), .IN3(\R[6][16] ), .IN2(\R[5][16] ), .IN4(
        \R[7][16] ), .S0(N190), .S1(n4084), .Q(n4051) );
  MUX21X1 U3124 ( .IN1(n4052), .IN2(n4051), .S(N191), .Q(N392) );
  MUX41X1 U3125 ( .IN1(\R[0][17] ), .IN3(\R[2][17] ), .IN2(\R[1][17] ), .IN4(
        \R[3][17] ), .S0(N190), .S1(n5715), .Q(n4054) );
  MUX21X1 U3126 ( .IN1(n4054), .IN2(n4053), .S(N191), .Q(N391) );
  MUX41X1 U3127 ( .IN1(\R[4][18] ), .IN3(\R[6][18] ), .IN2(\R[5][18] ), .IN4(
        \R[7][18] ), .S0(N190), .S1(n4086), .Q(n4055) );
  MUX21X1 U3128 ( .IN1(n4056), .IN2(n4055), .S(N191), .Q(N390) );
  MUX41X1 U3129 ( .IN1(\R[0][19] ), .IN3(\R[2][19] ), .IN2(\R[1][19] ), .IN4(
        \R[3][19] ), .S0(N190), .S1(n4083), .Q(n4058) );
  MUX21X1 U3130 ( .IN1(n4058), .IN2(n4057), .S(N191), .Q(N389) );
  MUX41X1 U3131 ( .IN1(\R[4][20] ), .IN3(\R[6][20] ), .IN2(\R[5][20] ), .IN4(
        \R[7][20] ), .S0(N190), .S1(n5715), .Q(n4059) );
  MUX21X1 U3132 ( .IN1(n4060), .IN2(n4059), .S(N191), .Q(N388) );
  MUX41X1 U3133 ( .IN1(\R[0][21] ), .IN3(\R[2][21] ), .IN2(\R[1][21] ), .IN4(
        \R[3][21] ), .S0(N190), .S1(n4085), .Q(n4062) );
  MUX21X1 U3134 ( .IN1(n4062), .IN2(n4061), .S(N191), .Q(N387) );
  MUX41X1 U3135 ( .IN1(\R[4][22] ), .IN3(\R[6][22] ), .IN2(\R[5][22] ), .IN4(
        \R[7][22] ), .S0(N190), .S1(n4083), .Q(n4063) );
  MUX21X1 U3136 ( .IN1(n4064), .IN2(n4063), .S(N191), .Q(N386) );
  MUX41X1 U3137 ( .IN1(\R[4][23] ), .IN3(\R[6][23] ), .IN2(\R[5][23] ), .IN4(
        \R[7][23] ), .S0(N190), .S1(n4083), .Q(n4065) );
  MUX41X1 U3138 ( .IN1(\R[0][23] ), .IN3(\R[2][23] ), .IN2(\R[1][23] ), .IN4(
        \R[3][23] ), .S0(N190), .S1(n4083), .Q(n4066) );
  MUX21X1 U3139 ( .IN1(n4066), .IN2(n4065), .S(N191), .Q(N385) );
  MUX21X1 U3140 ( .IN1(n4068), .IN2(n4067), .S(N191), .Q(N384) );
  MUX41X1 U3141 ( .IN1(\R[4][25] ), .IN3(\R[6][25] ), .IN2(\R[5][25] ), .IN4(
        \R[7][25] ), .S0(N190), .S1(n4084), .Q(n4069) );
  MUX41X1 U3142 ( .IN1(\R[0][25] ), .IN3(\R[2][25] ), .IN2(\R[1][25] ), .IN4(
        \R[3][25] ), .S0(N190), .S1(n4083), .Q(n4070) );
  MUX21X1 U3143 ( .IN1(n4070), .IN2(n4069), .S(N191), .Q(N383) );
  MUX41X1 U3144 ( .IN1(\R[0][26] ), .IN3(\R[2][26] ), .IN2(\R[1][26] ), .IN4(
        \R[3][26] ), .S0(N190), .S1(n4086), .Q(n4072) );
  MUX21X1 U3145 ( .IN1(n4072), .IN2(n4071), .S(N191), .Q(N382) );
  MUX41X1 U3146 ( .IN1(\R[4][27] ), .IN3(\R[6][27] ), .IN2(\R[5][27] ), .IN4(
        \R[7][27] ), .S0(N190), .S1(n4083), .Q(n4073) );
  MUX21X1 U3147 ( .IN1(n4074), .IN2(n4073), .S(N191), .Q(N381) );
  MUX41X1 U3148 ( .IN1(\R[0][28] ), .IN3(\R[2][28] ), .IN2(\R[1][28] ), .IN4(
        \R[3][28] ), .S0(N190), .S1(n4084), .Q(n4076) );
  MUX21X1 U3149 ( .IN1(n4076), .IN2(n4075), .S(N191), .Q(N380) );
  MUX41X1 U3150 ( .IN1(\R[4][29] ), .IN3(\R[6][29] ), .IN2(\R[5][29] ), .IN4(
        \R[7][29] ), .S0(N190), .S1(n4086), .Q(n4077) );
  MUX21X1 U3151 ( .IN1(n4078), .IN2(n4077), .S(N191), .Q(N379) );
  MUX41X1 U3152 ( .IN1(\R[0][30] ), .IN3(\R[2][30] ), .IN2(\R[1][30] ), .IN4(
        \R[3][30] ), .S0(N190), .S1(n4085), .Q(n4080) );
  MUX21X1 U3153 ( .IN1(n4080), .IN2(n4079), .S(N191), .Q(N378) );
  MUX41X1 U3154 ( .IN1(\R[4][31] ), .IN3(\R[6][31] ), .IN2(\R[5][31] ), .IN4(
        \R[7][31] ), .S0(N190), .S1(n5715), .Q(n4081) );
  MUX21X1 U3155 ( .IN1(n4082), .IN2(n4081), .S(N191), .Q(N377) );
  MUX41X1 U3156 ( .IN1(\R[4][0] ), .IN3(\R[6][0] ), .IN2(\R[5][0] ), .IN4(
        \R[7][0] ), .S0(N193), .S1(n4160), .Q(n4087) );
  MUX41X1 U3157 ( .IN1(\R[0][0] ), .IN3(\R[2][0] ), .IN2(\R[1][0] ), .IN4(
        \R[3][0] ), .S0(N193), .S1(n4159), .Q(n4088) );
  MUX21X1 U3158 ( .IN1(n4088), .IN2(n4087), .S(n5719), .Q(N440) );
  MUX41X1 U3159 ( .IN1(\R[4][1] ), .IN3(\R[6][1] ), .IN2(\R[5][1] ), .IN4(
        \R[7][1] ), .S0(N193), .S1(n4158), .Q(n4089) );
  MUX41X1 U3160 ( .IN1(\R[0][1] ), .IN3(\R[2][1] ), .IN2(\R[1][1] ), .IN4(
        \R[3][1] ), .S0(N193), .S1(n4157), .Q(n4090) );
  MUX21X1 U3161 ( .IN1(n4090), .IN2(n4089), .S(n4234), .Q(N439) );
  MUX41X1 U3162 ( .IN1(\R[4][2] ), .IN3(\R[6][2] ), .IN2(\R[5][2] ), .IN4(
        \R[7][2] ), .S0(N193), .S1(n4156), .Q(n4091) );
  MUX41X1 U3163 ( .IN1(\R[0][2] ), .IN3(\R[2][2] ), .IN2(\R[1][2] ), .IN4(
        \R[3][2] ), .S0(N193), .S1(n4155), .Q(n4092) );
  MUX21X1 U3164 ( .IN1(n4092), .IN2(n4091), .S(n4227), .Q(N438) );
  MUX41X1 U3165 ( .IN1(\R[4][3] ), .IN3(\R[6][3] ), .IN2(\R[5][3] ), .IN4(
        \R[7][3] ), .S0(N193), .S1(n4154), .Q(n4093) );
  MUX41X1 U3166 ( .IN1(\R[0][3] ), .IN3(\R[2][3] ), .IN2(\R[1][3] ), .IN4(
        \R[3][3] ), .S0(N193), .S1(n4153), .Q(n4094) );
  MUX21X1 U3167 ( .IN1(n4094), .IN2(n4093), .S(n4229), .Q(N437) );
  MUX41X1 U3168 ( .IN1(\R[4][4] ), .IN3(\R[6][4] ), .IN2(\R[5][4] ), .IN4(
        \R[7][4] ), .S0(N193), .S1(n4157), .Q(n4095) );
  MUX41X1 U3169 ( .IN1(\R[0][4] ), .IN3(\R[2][4] ), .IN2(\R[1][4] ), .IN4(
        \R[3][4] ), .S0(N193), .S1(n4152), .Q(n4096) );
  MUX21X1 U3170 ( .IN1(n4096), .IN2(n4095), .S(n4235), .Q(N436) );
  MUX41X1 U3171 ( .IN1(\R[4][5] ), .IN3(\R[6][5] ), .IN2(\R[5][5] ), .IN4(
        \R[7][5] ), .S0(N193), .S1(n4158), .Q(n4097) );
  MUX41X1 U3172 ( .IN1(\R[0][5] ), .IN3(\R[2][5] ), .IN2(\R[1][5] ), .IN4(
        \R[3][5] ), .S0(N193), .S1(n4153), .Q(n4098) );
  MUX21X1 U3173 ( .IN1(n4098), .IN2(n4097), .S(n4233), .Q(N435) );
  MUX41X1 U3174 ( .IN1(\R[4][6] ), .IN3(\R[6][6] ), .IN2(\R[5][6] ), .IN4(
        \R[7][6] ), .S0(N193), .S1(n5705), .Q(n4099) );
  MUX41X1 U3175 ( .IN1(\R[0][6] ), .IN3(\R[2][6] ), .IN2(\R[1][6] ), .IN4(
        \R[3][6] ), .S0(N193), .S1(n5705), .Q(n4100) );
  MUX21X1 U3176 ( .IN1(n4100), .IN2(n4099), .S(n4227), .Q(N434) );
  MUX41X1 U3177 ( .IN1(\R[4][7] ), .IN3(\R[6][7] ), .IN2(\R[5][7] ), .IN4(
        \R[7][7] ), .S0(N193), .S1(n4159), .Q(n4101) );
  MUX41X1 U3178 ( .IN1(\R[0][7] ), .IN3(\R[2][7] ), .IN2(\R[1][7] ), .IN4(
        \R[3][7] ), .S0(N193), .S1(n4153), .Q(n4102) );
  MUX21X1 U3179 ( .IN1(n4102), .IN2(n4101), .S(n4226), .Q(N433) );
  MUX41X1 U3180 ( .IN1(\R[4][8] ), .IN3(\R[6][8] ), .IN2(\R[5][8] ), .IN4(
        \R[7][8] ), .S0(N193), .S1(n4155), .Q(n4103) );
  MUX41X1 U3181 ( .IN1(\R[0][8] ), .IN3(\R[2][8] ), .IN2(\R[1][8] ), .IN4(
        \R[3][8] ), .S0(N193), .S1(n4159), .Q(n4104) );
  MUX21X1 U3182 ( .IN1(n4104), .IN2(n4103), .S(n4226), .Q(N432) );
  MUX41X1 U3183 ( .IN1(\R[4][9] ), .IN3(\R[6][9] ), .IN2(\R[5][9] ), .IN4(
        \R[7][9] ), .S0(N193), .S1(n4160), .Q(n4105) );
  MUX41X1 U3184 ( .IN1(\R[0][9] ), .IN3(\R[2][9] ), .IN2(\R[1][9] ), .IN4(
        \R[3][9] ), .S0(N193), .S1(n4151), .Q(n4106) );
  MUX21X1 U3185 ( .IN1(n4106), .IN2(n4105), .S(n4229), .Q(N431) );
  MUX41X1 U3186 ( .IN1(\R[4][10] ), .IN3(\R[6][10] ), .IN2(\R[5][10] ), .IN4(
        \R[7][10] ), .S0(N193), .S1(n4156), .Q(n4107) );
  MUX41X1 U3187 ( .IN1(\R[0][10] ), .IN3(\R[2][10] ), .IN2(\R[1][10] ), .IN4(
        \R[3][10] ), .S0(N193), .S1(n4151), .Q(n4108) );
  MUX21X1 U3188 ( .IN1(n4108), .IN2(n4107), .S(n4236), .Q(N430) );
  MUX41X1 U3189 ( .IN1(\R[4][11] ), .IN3(\R[6][11] ), .IN2(\R[5][11] ), .IN4(
        \R[7][11] ), .S0(N193), .S1(n4152), .Q(n4109) );
  MUX41X1 U3190 ( .IN1(\R[0][11] ), .IN3(\R[2][11] ), .IN2(\R[1][11] ), .IN4(
        \R[3][11] ), .S0(N193), .S1(n4158), .Q(n4110) );
  MUX21X1 U3191 ( .IN1(n4110), .IN2(n4109), .S(n4232), .Q(N429) );
  MUX41X1 U3192 ( .IN1(\R[4][12] ), .IN3(\R[6][12] ), .IN2(\R[5][12] ), .IN4(
        \R[7][12] ), .S0(N193), .S1(n4158), .Q(n4111) );
  MUX41X1 U3193 ( .IN1(\R[0][12] ), .IN3(\R[2][12] ), .IN2(\R[1][12] ), .IN4(
        \R[3][12] ), .S0(N193), .S1(n4153), .Q(n4112) );
  MUX21X1 U3194 ( .IN1(n4112), .IN2(n4111), .S(n4229), .Q(N428) );
  MUX41X1 U3195 ( .IN1(\R[4][13] ), .IN3(\R[6][13] ), .IN2(\R[5][13] ), .IN4(
        \R[7][13] ), .S0(N193), .S1(n4151), .Q(n4113) );
  MUX41X1 U3196 ( .IN1(\R[0][13] ), .IN3(\R[2][13] ), .IN2(\R[1][13] ), .IN4(
        \R[3][13] ), .S0(N193), .S1(n4159), .Q(n4114) );
  MUX21X1 U3197 ( .IN1(n4114), .IN2(n4113), .S(n4228), .Q(N427) );
  MUX41X1 U3198 ( .IN1(\R[4][14] ), .IN3(\R[6][14] ), .IN2(\R[5][14] ), .IN4(
        \R[7][14] ), .S0(N193), .S1(n4159), .Q(n4115) );
  MUX41X1 U3199 ( .IN1(\R[0][14] ), .IN3(\R[2][14] ), .IN2(\R[1][14] ), .IN4(
        \R[3][14] ), .S0(N193), .S1(n4155), .Q(n4116) );
  MUX21X1 U3200 ( .IN1(n4116), .IN2(n4115), .S(n4232), .Q(N426) );
  MUX41X1 U3201 ( .IN1(\R[4][15] ), .IN3(\R[6][15] ), .IN2(\R[5][15] ), .IN4(
        \R[7][15] ), .S0(N193), .S1(n4152), .Q(n4117) );
  MUX41X1 U3202 ( .IN1(\R[0][15] ), .IN3(\R[2][15] ), .IN2(\R[1][15] ), .IN4(
        \R[3][15] ), .S0(N193), .S1(n4154), .Q(n4118) );
  MUX21X1 U3203 ( .IN1(n4118), .IN2(n4117), .S(n4231), .Q(N425) );
  MUX41X1 U3204 ( .IN1(\R[4][16] ), .IN3(\R[6][16] ), .IN2(\R[5][16] ), .IN4(
        \R[7][16] ), .S0(N193), .S1(n4153), .Q(n4119) );
  MUX41X1 U3205 ( .IN1(\R[0][16] ), .IN3(\R[2][16] ), .IN2(\R[1][16] ), .IN4(
        \R[3][16] ), .S0(N193), .S1(n4154), .Q(n4120) );
  MUX21X1 U3206 ( .IN1(n4120), .IN2(n4119), .S(n4234), .Q(N424) );
  MUX41X1 U3207 ( .IN1(\R[4][17] ), .IN3(\R[6][17] ), .IN2(\R[5][17] ), .IN4(
        \R[7][17] ), .S0(N193), .S1(n4155), .Q(n4121) );
  MUX41X1 U3208 ( .IN1(\R[0][17] ), .IN3(\R[2][17] ), .IN2(\R[1][17] ), .IN4(
        \R[3][17] ), .S0(N193), .S1(n4156), .Q(n4122) );
  MUX21X1 U3209 ( .IN1(n4122), .IN2(n4121), .S(n4233), .Q(N423) );
  MUX41X1 U3210 ( .IN1(\R[4][18] ), .IN3(\R[6][18] ), .IN2(\R[5][18] ), .IN4(
        \R[7][18] ), .S0(N193), .S1(n4157), .Q(n4123) );
  MUX41X1 U3211 ( .IN1(\R[0][18] ), .IN3(\R[2][18] ), .IN2(\R[1][18] ), .IN4(
        \R[3][18] ), .S0(N193), .S1(n4158), .Q(n4124) );
  MUX21X1 U3212 ( .IN1(n4124), .IN2(n4123), .S(n4234), .Q(N422) );
  MUX41X1 U3213 ( .IN1(\R[4][19] ), .IN3(\R[6][19] ), .IN2(\R[5][19] ), .IN4(
        \R[7][19] ), .S0(N193), .S1(n4159), .Q(n4125) );
  MUX41X1 U3214 ( .IN1(\R[0][19] ), .IN3(\R[2][19] ), .IN2(\R[1][19] ), .IN4(
        \R[3][19] ), .S0(N193), .S1(n4160), .Q(n4126) );
  MUX21X1 U3215 ( .IN1(n4126), .IN2(n4125), .S(n4233), .Q(N421) );
  MUX41X1 U3216 ( .IN1(\R[4][20] ), .IN3(\R[6][20] ), .IN2(\R[5][20] ), .IN4(
        \R[7][20] ), .S0(N193), .S1(n4152), .Q(n4127) );
  MUX41X1 U3217 ( .IN1(\R[0][20] ), .IN3(\R[2][20] ), .IN2(\R[1][20] ), .IN4(
        \R[3][20] ), .S0(N193), .S1(n5705), .Q(n4128) );
  MUX21X1 U3218 ( .IN1(n4128), .IN2(n4127), .S(n4236), .Q(N420) );
  MUX41X1 U3219 ( .IN1(\R[4][21] ), .IN3(\R[6][21] ), .IN2(\R[5][21] ), .IN4(
        \R[7][21] ), .S0(N193), .S1(n5705), .Q(n4129) );
  MUX41X1 U3220 ( .IN1(\R[0][21] ), .IN3(\R[2][21] ), .IN2(\R[1][21] ), .IN4(
        \R[3][21] ), .S0(N193), .S1(n4152), .Q(n4130) );
  MUX21X1 U3221 ( .IN1(n4130), .IN2(n4129), .S(n4235), .Q(N419) );
  MUX41X1 U3222 ( .IN1(\R[4][22] ), .IN3(\R[6][22] ), .IN2(\R[5][22] ), .IN4(
        \R[7][22] ), .S0(N193), .S1(n4156), .Q(n4131) );
  MUX41X1 U3223 ( .IN1(\R[0][22] ), .IN3(\R[2][22] ), .IN2(\R[1][22] ), .IN4(
        \R[3][22] ), .S0(N193), .S1(n4157), .Q(n4132) );
  MUX21X1 U3224 ( .IN1(n4132), .IN2(n4131), .S(n4238), .Q(N418) );
  MUX41X1 U3225 ( .IN1(\R[4][23] ), .IN3(\R[6][23] ), .IN2(\R[5][23] ), .IN4(
        \R[7][23] ), .S0(N193), .S1(n4155), .Q(n4133) );
  MUX41X1 U3226 ( .IN1(\R[0][23] ), .IN3(\R[2][23] ), .IN2(\R[1][23] ), .IN4(
        \R[3][23] ), .S0(N193), .S1(n4151), .Q(n4134) );
  MUX21X1 U3227 ( .IN1(n4134), .IN2(n4133), .S(n4237), .Q(N417) );
  MUX41X1 U3228 ( .IN1(\R[4][24] ), .IN3(\R[6][24] ), .IN2(\R[5][24] ), .IN4(
        \R[7][24] ), .S0(N193), .S1(n4151), .Q(n4135) );
  MUX41X1 U3229 ( .IN1(\R[0][24] ), .IN3(\R[2][24] ), .IN2(\R[1][24] ), .IN4(
        \R[3][24] ), .S0(N193), .S1(n4160), .Q(n4136) );
  MUX21X1 U3230 ( .IN1(n4136), .IN2(n4135), .S(n4226), .Q(N416) );
  MUX41X1 U3231 ( .IN1(\R[4][25] ), .IN3(\R[6][25] ), .IN2(\R[5][25] ), .IN4(
        \R[7][25] ), .S0(N193), .S1(n4160), .Q(n4137) );
  MUX41X1 U3232 ( .IN1(\R[0][25] ), .IN3(\R[2][25] ), .IN2(\R[1][25] ), .IN4(
        \R[3][25] ), .S0(N193), .S1(n4157), .Q(n4138) );
  MUX21X1 U3233 ( .IN1(n4138), .IN2(n4137), .S(n4232), .Q(N415) );
  MUX41X1 U3234 ( .IN1(\R[4][26] ), .IN3(\R[6][26] ), .IN2(\R[5][26] ), .IN4(
        \R[7][26] ), .S0(N193), .S1(n4154), .Q(n4139) );
  MUX41X1 U3235 ( .IN1(\R[0][26] ), .IN3(\R[2][26] ), .IN2(\R[1][26] ), .IN4(
        \R[3][26] ), .S0(N193), .S1(n4155), .Q(n4140) );
  MUX21X1 U3236 ( .IN1(n4140), .IN2(n4139), .S(n4230), .Q(N414) );
  MUX41X1 U3237 ( .IN1(\R[4][27] ), .IN3(\R[6][27] ), .IN2(\R[5][27] ), .IN4(
        \R[7][27] ), .S0(N193), .S1(n4152), .Q(n4141) );
  MUX41X1 U3238 ( .IN1(\R[0][27] ), .IN3(\R[2][27] ), .IN2(\R[1][27] ), .IN4(
        \R[3][27] ), .S0(N193), .S1(n4156), .Q(n4142) );
  MUX21X1 U3239 ( .IN1(n4142), .IN2(n4141), .S(n5719), .Q(N413) );
  MUX41X1 U3240 ( .IN1(\R[4][28] ), .IN3(\R[6][28] ), .IN2(\R[5][28] ), .IN4(
        \R[7][28] ), .S0(N193), .S1(n4158), .Q(n4143) );
  MUX41X1 U3241 ( .IN1(\R[0][28] ), .IN3(\R[2][28] ), .IN2(\R[1][28] ), .IN4(
        \R[3][28] ), .S0(N193), .S1(n4154), .Q(n4144) );
  MUX21X1 U3242 ( .IN1(n4144), .IN2(n4143), .S(n4235), .Q(N412) );
  MUX41X1 U3243 ( .IN1(\R[4][29] ), .IN3(\R[6][29] ), .IN2(\R[5][29] ), .IN4(
        \R[7][29] ), .S0(N193), .S1(n4151), .Q(n4145) );
  MUX41X1 U3244 ( .IN1(\R[0][29] ), .IN3(\R[2][29] ), .IN2(\R[1][29] ), .IN4(
        \R[3][29] ), .S0(N193), .S1(n4156), .Q(n4146) );
  MUX21X1 U3245 ( .IN1(n4146), .IN2(n4145), .S(n4236), .Q(N411) );
  MUX41X1 U3246 ( .IN1(\R[4][30] ), .IN3(\R[6][30] ), .IN2(\R[5][30] ), .IN4(
        \R[7][30] ), .S0(N193), .S1(n4157), .Q(n4147) );
  MUX41X1 U3247 ( .IN1(\R[0][30] ), .IN3(\R[2][30] ), .IN2(\R[1][30] ), .IN4(
        \R[3][30] ), .S0(N193), .S1(n4153), .Q(n4148) );
  MUX21X1 U3248 ( .IN1(n4148), .IN2(n4147), .S(n4227), .Q(N410) );
  MUX41X1 U3249 ( .IN1(\R[4][31] ), .IN3(\R[6][31] ), .IN2(\R[5][31] ), .IN4(
        \R[7][31] ), .S0(N193), .S1(n4154), .Q(n4149) );
  MUX41X1 U3250 ( .IN1(\R[0][31] ), .IN3(\R[2][31] ), .IN2(\R[1][31] ), .IN4(
        \R[3][31] ), .S0(N193), .S1(n4160), .Q(n4150) );
  MUX21X1 U3251 ( .IN1(n4150), .IN2(n4149), .S(n4225), .Q(N409) );
  MUX41X1 U3252 ( .IN1(\R[4][0] ), .IN3(\R[6][0] ), .IN2(\R[5][0] ), .IN4(
        \R[7][0] ), .S0(N195), .S1(n4238), .Q(n4161) );
  MUX41X1 U3253 ( .IN1(\R[0][0] ), .IN3(\R[2][0] ), .IN2(\R[1][0] ), .IN4(
        \R[3][0] ), .S0(N195), .S1(n4233), .Q(n4162) );
  MUX21X1 U3254 ( .IN1(n4162), .IN2(n4161), .S(N196), .Q(N472) );
  MUX41X1 U3255 ( .IN1(\R[4][1] ), .IN3(\R[6][1] ), .IN2(\R[5][1] ), .IN4(
        \R[7][1] ), .S0(N195), .S1(n4237), .Q(n4163) );
  MUX41X1 U3256 ( .IN1(\R[0][1] ), .IN3(\R[2][1] ), .IN2(\R[1][1] ), .IN4(
        \R[3][1] ), .S0(N195), .S1(n4235), .Q(n4164) );
  MUX21X1 U3257 ( .IN1(n4164), .IN2(n4163), .S(N196), .Q(N471) );
  MUX41X1 U3258 ( .IN1(\R[4][2] ), .IN3(\R[6][2] ), .IN2(\R[5][2] ), .IN4(
        \R[7][2] ), .S0(N195), .S1(n4236), .Q(n4165) );
  MUX41X1 U3259 ( .IN1(\R[0][2] ), .IN3(\R[2][2] ), .IN2(\R[1][2] ), .IN4(
        \R[3][2] ), .S0(N195), .S1(n4237), .Q(n4166) );
  MUX21X1 U3260 ( .IN1(n4166), .IN2(n4165), .S(N196), .Q(N470) );
  MUX41X1 U3261 ( .IN1(\R[4][3] ), .IN3(\R[6][3] ), .IN2(\R[5][3] ), .IN4(
        \R[7][3] ), .S0(N195), .S1(n4235), .Q(n4167) );
  MUX41X1 U3262 ( .IN1(\R[0][3] ), .IN3(\R[2][3] ), .IN2(\R[1][3] ), .IN4(
        \R[3][3] ), .S0(N195), .S1(n4228), .Q(n4168) );
  MUX21X1 U3263 ( .IN1(n4168), .IN2(n4167), .S(N196), .Q(N469) );
  MUX41X1 U3264 ( .IN1(\R[4][4] ), .IN3(\R[6][4] ), .IN2(\R[5][4] ), .IN4(
        \R[7][4] ), .S0(N195), .S1(n4234), .Q(n4169) );
  MUX41X1 U3265 ( .IN1(\R[0][4] ), .IN3(\R[2][4] ), .IN2(\R[1][4] ), .IN4(
        \R[3][4] ), .S0(N195), .S1(n4228), .Q(n4170) );
  MUX21X1 U3266 ( .IN1(n4170), .IN2(n4169), .S(N196), .Q(N468) );
  MUX41X1 U3267 ( .IN1(\R[4][5] ), .IN3(\R[6][5] ), .IN2(\R[5][5] ), .IN4(
        \R[7][5] ), .S0(N195), .S1(n4233), .Q(n4171) );
  MUX41X1 U3268 ( .IN1(\R[0][5] ), .IN3(\R[2][5] ), .IN2(\R[1][5] ), .IN4(
        \R[3][5] ), .S0(N195), .S1(n4225), .Q(n4172) );
  MUX21X1 U3269 ( .IN1(n4172), .IN2(n4171), .S(N196), .Q(N467) );
  MUX41X1 U3270 ( .IN1(\R[4][6] ), .IN3(\R[6][6] ), .IN2(\R[5][6] ), .IN4(
        \R[7][6] ), .S0(N195), .S1(n4232), .Q(n4173) );
  MUX41X1 U3271 ( .IN1(\R[0][6] ), .IN3(\R[2][6] ), .IN2(\R[1][6] ), .IN4(
        \R[3][6] ), .S0(N195), .S1(n4227), .Q(n4174) );
  MUX21X1 U3272 ( .IN1(n4174), .IN2(n4173), .S(N196), .Q(N466) );
  MUX41X1 U3273 ( .IN1(\R[4][7] ), .IN3(\R[6][7] ), .IN2(\R[5][7] ), .IN4(
        \R[7][7] ), .S0(N195), .S1(n4231), .Q(n4175) );
  MUX41X1 U3274 ( .IN1(\R[0][7] ), .IN3(\R[2][7] ), .IN2(\R[1][7] ), .IN4(
        \R[3][7] ), .S0(N195), .S1(n4230), .Q(n4176) );
  MUX21X1 U3275 ( .IN1(n4176), .IN2(n4175), .S(N196), .Q(N465) );
  MUX41X1 U3276 ( .IN1(\R[4][8] ), .IN3(\R[6][8] ), .IN2(\R[5][8] ), .IN4(
        \R[7][8] ), .S0(N195), .S1(n4230), .Q(n4177) );
  MUX41X1 U3277 ( .IN1(\R[0][8] ), .IN3(\R[2][8] ), .IN2(\R[1][8] ), .IN4(
        \R[3][8] ), .S0(N195), .S1(n4232), .Q(n4178) );
  MUX21X1 U3278 ( .IN1(n4178), .IN2(n4177), .S(N196), .Q(N464) );
  MUX41X1 U3279 ( .IN1(\R[4][9] ), .IN3(\R[6][9] ), .IN2(\R[5][9] ), .IN4(
        \R[7][9] ), .S0(N195), .S1(n4229), .Q(n4179) );
  MUX41X1 U3280 ( .IN1(\R[0][9] ), .IN3(\R[2][9] ), .IN2(\R[1][9] ), .IN4(
        \R[3][9] ), .S0(N195), .S1(n4230), .Q(n4180) );
  MUX21X1 U3281 ( .IN1(n4180), .IN2(n4179), .S(N196), .Q(N463) );
  MUX41X1 U3282 ( .IN1(\R[4][10] ), .IN3(\R[6][10] ), .IN2(\R[5][10] ), .IN4(
        \R[7][10] ), .S0(N195), .S1(n4228), .Q(n4181) );
  MUX41X1 U3283 ( .IN1(\R[0][10] ), .IN3(\R[2][10] ), .IN2(\R[1][10] ), .IN4(
        \R[3][10] ), .S0(N195), .S1(n4228), .Q(n4182) );
  MUX21X1 U3284 ( .IN1(n4182), .IN2(n4181), .S(N196), .Q(N462) );
  MUX41X1 U3285 ( .IN1(\R[4][11] ), .IN3(\R[6][11] ), .IN2(\R[5][11] ), .IN4(
        \R[7][11] ), .S0(N195), .S1(n4238), .Q(n4183) );
  MUX41X1 U3286 ( .IN1(\R[0][11] ), .IN3(\R[2][11] ), .IN2(\R[1][11] ), .IN4(
        \R[3][11] ), .S0(N195), .S1(n4230), .Q(n4184) );
  MUX21X1 U3287 ( .IN1(n4184), .IN2(n4183), .S(N196), .Q(N461) );
  MUX41X1 U3288 ( .IN1(\R[4][12] ), .IN3(\R[6][12] ), .IN2(\R[5][12] ), .IN4(
        \R[7][12] ), .S0(N195), .S1(n4231), .Q(n4185) );
  MUX41X1 U3289 ( .IN1(\R[0][12] ), .IN3(\R[2][12] ), .IN2(\R[1][12] ), .IN4(
        \R[3][12] ), .S0(N195), .S1(n4232), .Q(n4186) );
  MUX21X1 U3290 ( .IN1(n4186), .IN2(n4185), .S(N196), .Q(N460) );
  MUX41X1 U3291 ( .IN1(\R[4][13] ), .IN3(\R[6][13] ), .IN2(\R[5][13] ), .IN4(
        \R[7][13] ), .S0(N195), .S1(n4234), .Q(n4187) );
  MUX41X1 U3292 ( .IN1(\R[0][13] ), .IN3(\R[2][13] ), .IN2(\R[1][13] ), .IN4(
        \R[3][13] ), .S0(N195), .S1(n4231), .Q(n4188) );
  MUX21X1 U3293 ( .IN1(n4188), .IN2(n4187), .S(N196), .Q(N459) );
  MUX41X1 U3294 ( .IN1(\R[4][14] ), .IN3(\R[6][14] ), .IN2(\R[5][14] ), .IN4(
        \R[7][14] ), .S0(N195), .S1(n4233), .Q(n4189) );
  MUX41X1 U3295 ( .IN1(\R[0][14] ), .IN3(\R[2][14] ), .IN2(\R[1][14] ), .IN4(
        \R[3][14] ), .S0(N195), .S1(n4227), .Q(n4190) );
  MUX21X1 U3296 ( .IN1(n4190), .IN2(n4189), .S(N196), .Q(N458) );
  MUX41X1 U3297 ( .IN1(\R[4][15] ), .IN3(\R[6][15] ), .IN2(\R[5][15] ), .IN4(
        \R[7][15] ), .S0(N195), .S1(n4237), .Q(n4191) );
  MUX41X1 U3298 ( .IN1(\R[0][15] ), .IN3(\R[2][15] ), .IN2(\R[1][15] ), .IN4(
        \R[3][15] ), .S0(N195), .S1(n4225), .Q(n4192) );
  MUX21X1 U3299 ( .IN1(n4192), .IN2(n4191), .S(N196), .Q(N457) );
  MUX41X1 U3300 ( .IN1(\R[4][16] ), .IN3(\R[6][16] ), .IN2(\R[5][16] ), .IN4(
        \R[7][16] ), .S0(N195), .S1(n4231), .Q(n4193) );
  MUX41X1 U3301 ( .IN1(\R[0][16] ), .IN3(\R[2][16] ), .IN2(\R[1][16] ), .IN4(
        \R[3][16] ), .S0(N195), .S1(n4226), .Q(n4194) );
  MUX21X1 U3302 ( .IN1(n4194), .IN2(n4193), .S(N196), .Q(N456) );
  MUX41X1 U3303 ( .IN1(\R[4][17] ), .IN3(\R[6][17] ), .IN2(\R[5][17] ), .IN4(
        \R[7][17] ), .S0(N195), .S1(n4236), .Q(n4195) );
  MUX41X1 U3304 ( .IN1(\R[0][17] ), .IN3(\R[2][17] ), .IN2(\R[1][17] ), .IN4(
        \R[3][17] ), .S0(N195), .S1(n4225), .Q(n4196) );
  MUX21X1 U3305 ( .IN1(n4196), .IN2(n4195), .S(N196), .Q(N455) );
  MUX41X1 U3306 ( .IN1(\R[4][18] ), .IN3(\R[6][18] ), .IN2(\R[5][18] ), .IN4(
        \R[7][18] ), .S0(N195), .S1(n4227), .Q(n4197) );
  MUX41X1 U3307 ( .IN1(\R[0][18] ), .IN3(\R[2][18] ), .IN2(\R[1][18] ), .IN4(
        \R[3][18] ), .S0(N195), .S1(n4236), .Q(n4198) );
  MUX21X1 U3308 ( .IN1(n4198), .IN2(n4197), .S(N196), .Q(N454) );
  MUX41X1 U3309 ( .IN1(\R[4][19] ), .IN3(\R[6][19] ), .IN2(\R[5][19] ), .IN4(
        \R[7][19] ), .S0(N195), .S1(n4226), .Q(n4199) );
  MUX41X1 U3310 ( .IN1(\R[0][19] ), .IN3(\R[2][19] ), .IN2(\R[1][19] ), .IN4(
        \R[3][19] ), .S0(N195), .S1(n4227), .Q(n4200) );
  MUX21X1 U3311 ( .IN1(n4200), .IN2(n4199), .S(N196), .Q(N453) );
  MUX41X1 U3312 ( .IN1(\R[4][20] ), .IN3(\R[6][20] ), .IN2(\R[5][20] ), .IN4(
        \R[7][20] ), .S0(N195), .S1(n4225), .Q(n4201) );
  MUX41X1 U3313 ( .IN1(\R[0][20] ), .IN3(\R[2][20] ), .IN2(\R[1][20] ), .IN4(
        \R[3][20] ), .S0(N195), .S1(n4235), .Q(n4202) );
  MUX21X1 U3314 ( .IN1(n4202), .IN2(n4201), .S(N196), .Q(N452) );
  MUX41X1 U3315 ( .IN1(\R[4][21] ), .IN3(\R[6][21] ), .IN2(\R[5][21] ), .IN4(
        \R[7][21] ), .S0(N195), .S1(n4238), .Q(n4203) );
  MUX41X1 U3316 ( .IN1(\R[0][21] ), .IN3(\R[2][21] ), .IN2(\R[1][21] ), .IN4(
        \R[3][21] ), .S0(N195), .S1(n4225), .Q(n4204) );
  MUX21X1 U3317 ( .IN1(n4204), .IN2(n4203), .S(N196), .Q(N451) );
  MUX41X1 U3318 ( .IN1(\R[4][22] ), .IN3(\R[6][22] ), .IN2(\R[5][22] ), .IN4(
        \R[7][22] ), .S0(N195), .S1(n4229), .Q(n4205) );
  MUX41X1 U3319 ( .IN1(\R[0][22] ), .IN3(\R[2][22] ), .IN2(\R[1][22] ), .IN4(
        \R[3][22] ), .S0(N195), .S1(n4230), .Q(n4206) );
  MUX21X1 U3320 ( .IN1(n4206), .IN2(n4205), .S(N196), .Q(N450) );
  MUX41X1 U3321 ( .IN1(\R[4][23] ), .IN3(\R[6][23] ), .IN2(\R[5][23] ), .IN4(
        \R[7][23] ), .S0(N195), .S1(n4226), .Q(n4207) );
  MUX41X1 U3322 ( .IN1(\R[0][23] ), .IN3(\R[2][23] ), .IN2(\R[1][23] ), .IN4(
        \R[3][23] ), .S0(N195), .S1(n4229), .Q(n4208) );
  MUX21X1 U3323 ( .IN1(n4208), .IN2(n4207), .S(N196), .Q(N449) );
  MUX41X1 U3324 ( .IN1(\R[4][24] ), .IN3(\R[6][24] ), .IN2(\R[5][24] ), .IN4(
        \R[7][24] ), .S0(N195), .S1(n5719), .Q(n4209) );
  MUX41X1 U3325 ( .IN1(\R[0][24] ), .IN3(\R[2][24] ), .IN2(\R[1][24] ), .IN4(
        \R[3][24] ), .S0(N195), .S1(n4235), .Q(n4210) );
  MUX21X1 U3326 ( .IN1(n4210), .IN2(n4209), .S(N196), .Q(N448) );
  MUX41X1 U3327 ( .IN1(\R[4][25] ), .IN3(\R[6][25] ), .IN2(\R[5][25] ), .IN4(
        \R[7][25] ), .S0(N195), .S1(n4226), .Q(n4211) );
  MUX41X1 U3328 ( .IN1(\R[0][25] ), .IN3(\R[2][25] ), .IN2(\R[1][25] ), .IN4(
        \R[3][25] ), .S0(N195), .S1(n4228), .Q(n4212) );
  MUX21X1 U3329 ( .IN1(n4212), .IN2(n4211), .S(N196), .Q(N447) );
  MUX41X1 U3330 ( .IN1(\R[4][26] ), .IN3(\R[6][26] ), .IN2(\R[5][26] ), .IN4(
        \R[7][26] ), .S0(N195), .S1(n4231), .Q(n4213) );
  MUX41X1 U3331 ( .IN1(\R[0][26] ), .IN3(\R[2][26] ), .IN2(\R[1][26] ), .IN4(
        \R[3][26] ), .S0(N195), .S1(n4238), .Q(n4214) );
  MUX21X1 U3332 ( .IN1(n4214), .IN2(n4213), .S(N196), .Q(N446) );
  MUX41X1 U3333 ( .IN1(\R[4][27] ), .IN3(\R[6][27] ), .IN2(\R[5][27] ), .IN4(
        \R[7][27] ), .S0(N195), .S1(n4237), .Q(n4215) );
  MUX41X1 U3334 ( .IN1(\R[0][27] ), .IN3(\R[2][27] ), .IN2(\R[1][27] ), .IN4(
        \R[3][27] ), .S0(N195), .S1(n4236), .Q(n4216) );
  MUX21X1 U3335 ( .IN1(n4216), .IN2(n4215), .S(N196), .Q(N445) );
  MUX41X1 U3336 ( .IN1(\R[4][28] ), .IN3(\R[6][28] ), .IN2(\R[5][28] ), .IN4(
        \R[7][28] ), .S0(N195), .S1(n4229), .Q(n4217) );
  MUX41X1 U3337 ( .IN1(\R[0][28] ), .IN3(\R[2][28] ), .IN2(\R[1][28] ), .IN4(
        \R[3][28] ), .S0(N195), .S1(n4234), .Q(n4218) );
  MUX21X1 U3338 ( .IN1(n4218), .IN2(n4217), .S(N196), .Q(N444) );
  MUX41X1 U3339 ( .IN1(\R[4][29] ), .IN3(\R[6][29] ), .IN2(\R[5][29] ), .IN4(
        \R[7][29] ), .S0(N195), .S1(n4237), .Q(n4219) );
  MUX41X1 U3340 ( .IN1(\R[0][29] ), .IN3(\R[2][29] ), .IN2(\R[1][29] ), .IN4(
        \R[3][29] ), .S0(N195), .S1(n4234), .Q(n4220) );
  MUX21X1 U3341 ( .IN1(n4220), .IN2(n4219), .S(N196), .Q(N443) );
  MUX41X1 U3342 ( .IN1(\R[4][30] ), .IN3(\R[6][30] ), .IN2(\R[5][30] ), .IN4(
        \R[7][30] ), .S0(N195), .S1(n5719), .Q(n4221) );
  MUX41X1 U3343 ( .IN1(\R[0][30] ), .IN3(\R[2][30] ), .IN2(\R[1][30] ), .IN4(
        \R[3][30] ), .S0(N195), .S1(n4233), .Q(n4222) );
  MUX21X1 U3344 ( .IN1(n4222), .IN2(n4221), .S(N196), .Q(N442) );
  MUX41X1 U3345 ( .IN1(\R[4][31] ), .IN3(\R[6][31] ), .IN2(\R[5][31] ), .IN4(
        \R[7][31] ), .S0(N195), .S1(n4232), .Q(n4223) );
  MUX41X1 U3346 ( .IN1(\R[0][31] ), .IN3(\R[2][31] ), .IN2(\R[1][31] ), .IN4(
        \R[3][31] ), .S0(N195), .S1(n4238), .Q(n4224) );
  MUX21X1 U3347 ( .IN1(n4224), .IN2(n4223), .S(N196), .Q(N441) );
  OR2X1 U3348 ( .IN1(n4239), .IN2(n4240), .Q(n3791) );
  MUX21X1 U3349 ( .IN1(n4241), .IN2(instruction[9]), .S(reset_n), .Q(n4240) );
  OR2X1 U3350 ( .IN1(n4239), .IN2(n4242), .Q(n3790) );
  MUX21X1 U3351 ( .IN1(n4243), .IN2(instruction[10]), .S(reset_n), .Q(n4242)
         );
  OR2X1 U3352 ( .IN1(n4239), .IN2(n4244), .Q(n3789) );
  MUX21X1 U3353 ( .IN1(n4245), .IN2(instruction[11]), .S(reset_n), .Q(n4244)
         );
  OR2X1 U3354 ( .IN1(n4239), .IN2(n4246), .Q(n3788) );
  MUX21X1 U3355 ( .IN1(IF_IR[12]), .IN2(instruction[12]), .S(reset_n), .Q(
        n4246) );
  OR2X1 U3356 ( .IN1(n4239), .IN2(n4247), .Q(n3787) );
  MUX21X1 U3357 ( .IN1(n4248), .IN2(instruction[14]), .S(reset_n), .Q(n4247)
         );
  OR2X1 U3358 ( .IN1(n4239), .IN2(n4249), .Q(n3786) );
  MUX21X1 U3359 ( .IN1(n4250), .IN2(instruction[15]), .S(reset_n), .Q(n4249)
         );
  INVX0 U3360 ( .INP(n4251), .ZN(n4239) );
  AO22X1 U3361 ( .IN1(n4252), .IN2(n4253), .IN3(instruction[13]), .IN4(n4254), 
        .Q(n3785) );
  MUX21X1 U3362 ( .IN1(N376), .IN2(ID_Rn[0]), .S(n4255), .Q(n3784) );
  MUX21X1 U3363 ( .IN1(N375), .IN2(ID_Rn[1]), .S(n4255), .Q(n3783) );
  MUX21X1 U3364 ( .IN1(N374), .IN2(ID_Rn[2]), .S(n4255), .Q(n3782) );
  MUX21X1 U3365 ( .IN1(N373), .IN2(ID_Rn[3]), .S(n4255), .Q(n3781) );
  MUX21X1 U3366 ( .IN1(N372), .IN2(ID_Rn[4]), .S(n4255), .Q(n3780) );
  MUX21X1 U3367 ( .IN1(N371), .IN2(ID_Rn[5]), .S(n4255), .Q(n3779) );
  MUX21X1 U3368 ( .IN1(N370), .IN2(ID_Rn[6]), .S(n4255), .Q(n3778) );
  MUX21X1 U3369 ( .IN1(N369), .IN2(ID_Rn[7]), .S(n4255), .Q(n3777) );
  MUX21X1 U3370 ( .IN1(N368), .IN2(ID_Rn[8]), .S(n4255), .Q(n3776) );
  MUX21X1 U3371 ( .IN1(N367), .IN2(ID_Rn[9]), .S(n4255), .Q(n3775) );
  MUX21X1 U3372 ( .IN1(N366), .IN2(ID_Rn[10]), .S(n4255), .Q(n3774) );
  MUX21X1 U3373 ( .IN1(N365), .IN2(ID_Rn[11]), .S(n4255), .Q(n3773) );
  MUX21X1 U3374 ( .IN1(N364), .IN2(ID_Rn[12]), .S(n4255), .Q(n3772) );
  MUX21X1 U3375 ( .IN1(N363), .IN2(ID_Rn[13]), .S(n4255), .Q(n3771) );
  MUX21X1 U3376 ( .IN1(N362), .IN2(ID_Rn[14]), .S(n4255), .Q(n3770) );
  MUX21X1 U3377 ( .IN1(N361), .IN2(ID_Rn[15]), .S(n4255), .Q(n3769) );
  MUX21X1 U3378 ( .IN1(N360), .IN2(ID_Rn[16]), .S(n4255), .Q(n3768) );
  MUX21X1 U3379 ( .IN1(N359), .IN2(ID_Rn[17]), .S(n4255), .Q(n3767) );
  MUX21X1 U3380 ( .IN1(N358), .IN2(ID_Rn[18]), .S(n4255), .Q(n3766) );
  MUX21X1 U3381 ( .IN1(N357), .IN2(ID_Rn[19]), .S(n4255), .Q(n3765) );
  MUX21X1 U3382 ( .IN1(N356), .IN2(ID_Rn[20]), .S(n4255), .Q(n3764) );
  MUX21X1 U3383 ( .IN1(N355), .IN2(ID_Rn[21]), .S(n4255), .Q(n3763) );
  MUX21X1 U3384 ( .IN1(N354), .IN2(ID_Rn[22]), .S(n4255), .Q(n3762) );
  MUX21X1 U3385 ( .IN1(N353), .IN2(ID_Rn[23]), .S(n4255), .Q(n3761) );
  MUX21X1 U3386 ( .IN1(N352), .IN2(ID_Rn[24]), .S(n4255), .Q(n3760) );
  MUX21X1 U3387 ( .IN1(N351), .IN2(ID_Rn[25]), .S(n4255), .Q(n3759) );
  MUX21X1 U3388 ( .IN1(N350), .IN2(ID_Rn[26]), .S(n4255), .Q(n3758) );
  MUX21X1 U3389 ( .IN1(N349), .IN2(ID_Rn[27]), .S(n4255), .Q(n3757) );
  MUX21X1 U3390 ( .IN1(N348), .IN2(ID_Rn[28]), .S(n4255), .Q(n3756) );
  MUX21X1 U3391 ( .IN1(N347), .IN2(ID_Rn[29]), .S(n4255), .Q(n3755) );
  MUX21X1 U3392 ( .IN1(N346), .IN2(ID_Rn[30]), .S(n4255), .Q(n3754) );
  MUX21X1 U3393 ( .IN1(N345), .IN2(ID_Rn[31]), .S(n4255), .Q(n3753) );
  AOI21X1 U3394 ( .IN1(n4256), .IN2(n3797), .IN3(n4257), .QN(n4255) );
  MUX21X1 U3395 ( .IN1(n3803), .IN2(N767), .S(n4258), .Q(n3752) );
  MUX21X1 U3396 ( .IN1(n3843), .IN2(N768), .S(n4258), .Q(n3751) );
  MUX21X1 U3397 ( .IN1(n3805), .IN2(N769), .S(n4258), .Q(n3750) );
  MUX21X1 U3398 ( .IN1(n3804), .IN2(N771), .S(n4258), .Q(n3749) );
  NAND2X0 U3399 ( .IN1(n4259), .IN2(n4251), .QN(n3748) );
  MUX21X1 U3400 ( .IN1(n5706), .IN2(n5722), .S(reset_n), .Q(n4259) );
  MUX21X1 U3401 ( .IN1(n3844), .IN2(N772), .S(n4258), .Q(n3747) );
  AO22X1 U3402 ( .IN1(n5719), .IN2(n4253), .IN3(instruction[8]), .IN4(n4254), 
        .Q(n3746) );
  AO22X1 U3403 ( .IN1(n4260), .IN2(n4253), .IN3(instruction[7]), .IN4(n4254), 
        .Q(n3745) );
  MUX21X1 U3404 ( .IN1(n4260), .IN2(ID_imm_offset[7]), .S(n4261), .Q(n3744) );
  AO22X1 U3405 ( .IN1(n5705), .IN2(n4253), .IN3(instruction[6]), .IN4(n4254), 
        .Q(n3743) );
  AO222X1 U3406 ( .IN1(N440), .IN2(n4262), .IN3(n4263), .IN4(N376), .IN5(n4264), .IN6(n4265), .Q(n3742) );
  AO222X1 U3407 ( .IN1(N439), .IN2(n4262), .IN3(n4263), .IN4(N375), .IN5(n4264), .IN6(n4266), .Q(n3741) );
  AO222X1 U3408 ( .IN1(N438), .IN2(n4262), .IN3(n4263), .IN4(N374), .IN5(n4264), .IN6(n4267), .Q(n3740) );
  AO222X1 U3409 ( .IN1(N437), .IN2(n4262), .IN3(n4263), .IN4(N373), .IN5(n4264), .IN6(n4268), .Q(n3739) );
  AO222X1 U3410 ( .IN1(N436), .IN2(n4262), .IN3(n4263), .IN4(N372), .IN5(n4264), .IN6(n4269), .Q(n3738) );
  AO222X1 U3411 ( .IN1(N435), .IN2(n4262), .IN3(n4263), .IN4(N371), .IN5(n4264), .IN6(n4270), .Q(n3737) );
  AO222X1 U3412 ( .IN1(N434), .IN2(n4262), .IN3(n4263), .IN4(N370), .IN5(n4264), .IN6(n4271), .Q(n3736) );
  AO222X1 U3413 ( .IN1(N433), .IN2(n4262), .IN3(n4263), .IN4(N369), .IN5(n4264), .IN6(n4272), .Q(n3735) );
  AO222X1 U3414 ( .IN1(N432), .IN2(n4262), .IN3(n4263), .IN4(N368), .IN5(n4264), .IN6(n4273), .Q(n3734) );
  AO222X1 U3415 ( .IN1(N431), .IN2(n4262), .IN3(n4263), .IN4(N367), .IN5(n4264), .IN6(n4274), .Q(n3733) );
  AO222X1 U3416 ( .IN1(N430), .IN2(n4262), .IN3(n4263), .IN4(N366), .IN5(n4264), .IN6(n4275), .Q(n3732) );
  AO222X1 U3417 ( .IN1(N429), .IN2(n4262), .IN3(n4263), .IN4(N365), .IN5(n4264), .IN6(n4276), .Q(n3731) );
  AO222X1 U3418 ( .IN1(N428), .IN2(n4262), .IN3(n4263), .IN4(N364), .IN5(n4264), .IN6(n4277), .Q(n3730) );
  AO222X1 U3419 ( .IN1(N427), .IN2(n4262), .IN3(n4263), .IN4(N363), .IN5(n4264), .IN6(n4278), .Q(n3729) );
  AO222X1 U3420 ( .IN1(N426), .IN2(n4262), .IN3(n4263), .IN4(N362), .IN5(n4264), .IN6(n4279), .Q(n3728) );
  AO222X1 U3421 ( .IN1(N425), .IN2(n4262), .IN3(n4263), .IN4(N361), .IN5(n4264), .IN6(n4280), .Q(n3727) );
  AO222X1 U3422 ( .IN1(N424), .IN2(n4262), .IN3(n4263), .IN4(N360), .IN5(n4264), .IN6(n4281), .Q(n3726) );
  AO222X1 U3423 ( .IN1(N423), .IN2(n4262), .IN3(n4263), .IN4(N359), .IN5(n4264), .IN6(n4282), .Q(n3725) );
  AO222X1 U3424 ( .IN1(N422), .IN2(n4262), .IN3(n4263), .IN4(N358), .IN5(n4264), .IN6(n4283), .Q(n3724) );
  AO222X1 U3425 ( .IN1(N421), .IN2(n4262), .IN3(n4263), .IN4(N357), .IN5(n4264), .IN6(n4284), .Q(n3723) );
  AO222X1 U3426 ( .IN1(N420), .IN2(n4262), .IN3(n4263), .IN4(N356), .IN5(n4264), .IN6(n4285), .Q(n3722) );
  AO222X1 U3427 ( .IN1(N419), .IN2(n4262), .IN3(n4263), .IN4(N355), .IN5(n4264), .IN6(n4286), .Q(n3721) );
  AO222X1 U3428 ( .IN1(N418), .IN2(n4262), .IN3(n4263), .IN4(N354), .IN5(n4264), .IN6(n4287), .Q(n3720) );
  AO222X1 U3429 ( .IN1(N417), .IN2(n4262), .IN3(n4263), .IN4(N353), .IN5(n4264), .IN6(n4288), .Q(n3719) );
  AO222X1 U3430 ( .IN1(N416), .IN2(n4262), .IN3(n4263), .IN4(N352), .IN5(n4264), .IN6(n4289), .Q(n3718) );
  AO222X1 U3431 ( .IN1(N415), .IN2(n4262), .IN3(n4263), .IN4(N351), .IN5(n4264), .IN6(n4290), .Q(n3717) );
  AO222X1 U3432 ( .IN1(N414), .IN2(n4262), .IN3(n4263), .IN4(N350), .IN5(n4264), .IN6(n4291), .Q(n3716) );
  AO222X1 U3433 ( .IN1(N413), .IN2(n4262), .IN3(n4263), .IN4(N349), .IN5(n4264), .IN6(n4292), .Q(n3715) );
  AO222X1 U3434 ( .IN1(N412), .IN2(n4262), .IN3(n4263), .IN4(N348), .IN5(n4264), .IN6(n4293), .Q(n3714) );
  AO222X1 U3435 ( .IN1(N411), .IN2(n4262), .IN3(n4263), .IN4(N347), .IN5(n4264), .IN6(n4294), .Q(n3713) );
  AO222X1 U3436 ( .IN1(N410), .IN2(n4262), .IN3(n4263), .IN4(N346), .IN5(n4264), .IN6(n4295), .Q(n3712) );
  AO222X1 U3437 ( .IN1(N409), .IN2(n4262), .IN3(n4263), .IN4(N345), .IN5(n4264), .IN6(n4296), .Q(n3711) );
  AND3X1 U3438 ( .IN1(n4297), .IN2(n5738), .IN3(n4298), .Q(n4263) );
  NAND2X0 U3439 ( .IN1(n4299), .IN2(n4248), .QN(n4297) );
  AND2X1 U3440 ( .IN1(n4257), .IN2(n4298), .Q(n4262) );
  INVX0 U3441 ( .INP(n4264), .ZN(n4298) );
  NAND3X0 U3442 ( .IN1(n4300), .IN2(n4301), .IN3(n4302), .QN(n4264) );
  NAND2X0 U3443 ( .IN1(N498), .IN2(n4243), .QN(n4301) );
  AOI21X1 U3444 ( .IN1(n4303), .IN2(n4304), .IN3(n4305), .QN(n4257) );
  MUX21X1 U3445 ( .IN1(n4306), .IN2(n5738), .S(n3132), .Q(n4303) );
  MUX21X1 U3446 ( .IN1(n3807), .IN2(n4307), .S(n4258), .Q(n3710) );
  AND2X1 U3447 ( .IN1(n4308), .IN2(n4309), .Q(n4258) );
  NAND4X0 U3448 ( .IN1(n3132), .IN2(N498), .IN3(n4252), .IN4(n4250), .QN(n4309) );
  MUX21X1 U3449 ( .IN1(n4310), .IN2(n4311), .S(n3797), .Q(n4308) );
  NAND2X0 U3450 ( .IN1(n4312), .IN2(n4250), .QN(n4311) );
  INVX0 U3451 ( .INP(n4256), .ZN(n4310) );
  AO221X1 U3452 ( .IN1(n4313), .IN2(n5739), .IN3(n3799), .IN4(n4314), .IN5(
        n4315), .Q(n4307) );
  AO22X1 U3453 ( .IN1(n4316), .IN2(n4248), .IN3(n4317), .IN4(N688), .Q(n4315)
         );
  NOR2X0 U3454 ( .IN1(n3131), .IN2(n3130), .QN(n4317) );
  NAND4X0 U3455 ( .IN1(n3131), .IN2(n4318), .IN3(n4319), .IN4(n4306), .QN(
        n4316) );
  INVX0 U3456 ( .INP(n4300), .ZN(n4313) );
  NAND2X0 U3457 ( .IN1(n4320), .IN2(n4248), .QN(n4300) );
  NAND2X0 U3458 ( .IN1(n4321), .IN2(n4251), .QN(n3709) );
  MUX21X1 U3459 ( .IN1(n5710), .IN2(n5720), .S(reset_n), .Q(n4321) );
  AO222X1 U3460 ( .IN1(N472), .IN2(n4322), .IN3(N408), .IN4(n4323), .IN5(n4324), .IN6(n4325), .Q(n3708) );
  MUX21X1 U3461 ( .IN1(n5740), .IN2(n4325), .S(n4326), .Q(n3707) );
  AO222X1 U3462 ( .IN1(N471), .IN2(n4322), .IN3(N407), .IN4(n4323), .IN5(n4324), .IN6(n4327), .Q(n3706) );
  MUX21X1 U3463 ( .IN1(n5741), .IN2(n4327), .S(n4326), .Q(n3705) );
  AO222X1 U3464 ( .IN1(N470), .IN2(n4322), .IN3(N406), .IN4(n4323), .IN5(n4324), .IN6(n4328), .Q(n3704) );
  MUX21X1 U3465 ( .IN1(n5742), .IN2(n4328), .S(n4326), .Q(n3703) );
  AO222X1 U3466 ( .IN1(N469), .IN2(n4322), .IN3(N405), .IN4(n4323), .IN5(n4324), .IN6(n4329), .Q(n3702) );
  MUX21X1 U3467 ( .IN1(n5743), .IN2(n4329), .S(n4326), .Q(n3701) );
  AO222X1 U3468 ( .IN1(N468), .IN2(n4322), .IN3(N404), .IN4(n4323), .IN5(n4324), .IN6(n4330), .Q(n3700) );
  MUX21X1 U3469 ( .IN1(n5744), .IN2(n4330), .S(n4326), .Q(n3699) );
  AO222X1 U3470 ( .IN1(N467), .IN2(n4322), .IN3(N403), .IN4(n4323), .IN5(n4324), .IN6(n4331), .Q(n3698) );
  MUX21X1 U3471 ( .IN1(n5745), .IN2(n4331), .S(n4326), .Q(n3697) );
  AO222X1 U3472 ( .IN1(N466), .IN2(n4322), .IN3(N402), .IN4(n4323), .IN5(n4324), .IN6(n4332), .Q(n3696) );
  MUX21X1 U3473 ( .IN1(n5746), .IN2(n4332), .S(n4326), .Q(n3695) );
  AO222X1 U3474 ( .IN1(N465), .IN2(n4322), .IN3(N401), .IN4(n4323), .IN5(n4324), .IN6(n4333), .Q(n3694) );
  MUX21X1 U3475 ( .IN1(n5747), .IN2(n4333), .S(n4326), .Q(n3693) );
  AO222X1 U3476 ( .IN1(N464), .IN2(n4322), .IN3(N400), .IN4(n4323), .IN5(n4324), .IN6(n4334), .Q(n3692) );
  MUX21X1 U3477 ( .IN1(n5748), .IN2(n4334), .S(n4326), .Q(n3691) );
  AO222X1 U3478 ( .IN1(N463), .IN2(n4322), .IN3(N399), .IN4(n4323), .IN5(n4324), .IN6(n4335), .Q(n3690) );
  MUX21X1 U3479 ( .IN1(n5749), .IN2(n4335), .S(n4326), .Q(n3689) );
  AO222X1 U3480 ( .IN1(N462), .IN2(n4322), .IN3(N398), .IN4(n4323), .IN5(n4324), .IN6(n4336), .Q(n3688) );
  MUX21X1 U3481 ( .IN1(n5750), .IN2(n4336), .S(n4326), .Q(n3687) );
  AO222X1 U3482 ( .IN1(N461), .IN2(n4322), .IN3(N397), .IN4(n4323), .IN5(n4324), .IN6(n4337), .Q(n3686) );
  MUX21X1 U3483 ( .IN1(n5751), .IN2(n4337), .S(n4326), .Q(n3685) );
  AO222X1 U3484 ( .IN1(N460), .IN2(n4322), .IN3(N396), .IN4(n4323), .IN5(n4324), .IN6(n4338), .Q(n3684) );
  MUX21X1 U3485 ( .IN1(n5752), .IN2(n4338), .S(n4326), .Q(n3683) );
  AO222X1 U3486 ( .IN1(N459), .IN2(n4322), .IN3(N395), .IN4(n4323), .IN5(n4324), .IN6(n4339), .Q(n3682) );
  MUX21X1 U3487 ( .IN1(n5753), .IN2(n4339), .S(n4326), .Q(n3681) );
  AO222X1 U3488 ( .IN1(N458), .IN2(n4322), .IN3(N394), .IN4(n4323), .IN5(n4324), .IN6(n4340), .Q(n3680) );
  MUX21X1 U3489 ( .IN1(n5754), .IN2(n4340), .S(n4326), .Q(n3679) );
  AO222X1 U3490 ( .IN1(N457), .IN2(n4322), .IN3(N393), .IN4(n4323), .IN5(n4324), .IN6(n4341), .Q(n3678) );
  MUX21X1 U3491 ( .IN1(n5755), .IN2(n4341), .S(n4326), .Q(n3677) );
  AO222X1 U3492 ( .IN1(N456), .IN2(n4322), .IN3(N392), .IN4(n4323), .IN5(n4324), .IN6(n4342), .Q(n3676) );
  MUX21X1 U3493 ( .IN1(n5756), .IN2(n4342), .S(n4326), .Q(n3675) );
  AO222X1 U3494 ( .IN1(N455), .IN2(n4322), .IN3(N391), .IN4(n4323), .IN5(n4324), .IN6(n4343), .Q(n3674) );
  MUX21X1 U3495 ( .IN1(n5757), .IN2(n4343), .S(n4326), .Q(n3673) );
  AO222X1 U3496 ( .IN1(N454), .IN2(n4322), .IN3(N390), .IN4(n4323), .IN5(n4324), .IN6(n4344), .Q(n3672) );
  MUX21X1 U3497 ( .IN1(n5758), .IN2(n4344), .S(n4326), .Q(n3671) );
  AO222X1 U3498 ( .IN1(N453), .IN2(n4322), .IN3(N389), .IN4(n4323), .IN5(n4324), .IN6(n4345), .Q(n3670) );
  MUX21X1 U3499 ( .IN1(n5759), .IN2(n4345), .S(n4326), .Q(n3669) );
  AO222X1 U3500 ( .IN1(N452), .IN2(n4322), .IN3(N388), .IN4(n4323), .IN5(n4324), .IN6(n4346), .Q(n3668) );
  MUX21X1 U3501 ( .IN1(n5760), .IN2(n4346), .S(n4326), .Q(n3667) );
  AO222X1 U3502 ( .IN1(N451), .IN2(n4322), .IN3(N387), .IN4(n4323), .IN5(n4324), .IN6(n4347), .Q(n3666) );
  MUX21X1 U3503 ( .IN1(n5761), .IN2(n4347), .S(n4326), .Q(n3665) );
  AO222X1 U3504 ( .IN1(N450), .IN2(n4322), .IN3(N386), .IN4(n4323), .IN5(n4324), .IN6(n4348), .Q(n3664) );
  MUX21X1 U3505 ( .IN1(n5762), .IN2(n4348), .S(n4326), .Q(n3663) );
  AO222X1 U3506 ( .IN1(N449), .IN2(n4322), .IN3(N385), .IN4(n4323), .IN5(n4324), .IN6(n4349), .Q(n3662) );
  MUX21X1 U3507 ( .IN1(n5763), .IN2(n4349), .S(n4326), .Q(n3661) );
  AO222X1 U3508 ( .IN1(N448), .IN2(n4322), .IN3(N384), .IN4(n4323), .IN5(n4324), .IN6(n4350), .Q(n3660) );
  MUX21X1 U3509 ( .IN1(n5764), .IN2(n4350), .S(n4326), .Q(n3659) );
  AO222X1 U3510 ( .IN1(N447), .IN2(n4322), .IN3(N383), .IN4(n4323), .IN5(n4324), .IN6(n4351), .Q(n3658) );
  MUX21X1 U3511 ( .IN1(n5765), .IN2(n4351), .S(n4326), .Q(n3657) );
  AO222X1 U3512 ( .IN1(N446), .IN2(n4322), .IN3(N382), .IN4(n4323), .IN5(n4324), .IN6(n4352), .Q(n3656) );
  MUX21X1 U3513 ( .IN1(n5766), .IN2(n4352), .S(n4326), .Q(n3655) );
  AO222X1 U3514 ( .IN1(N445), .IN2(n4322), .IN3(N381), .IN4(n4323), .IN5(n4324), .IN6(n4353), .Q(n3654) );
  MUX21X1 U3515 ( .IN1(n5767), .IN2(n4353), .S(n4326), .Q(n3653) );
  AO222X1 U3516 ( .IN1(N444), .IN2(n4322), .IN3(N380), .IN4(n4323), .IN5(n4324), .IN6(n4354), .Q(n3652) );
  MUX21X1 U3517 ( .IN1(n5768), .IN2(n4354), .S(n4326), .Q(n3651) );
  AO222X1 U3518 ( .IN1(N443), .IN2(n4322), .IN3(N379), .IN4(n4323), .IN5(n4324), .IN6(n4355), .Q(n3650) );
  MUX21X1 U3519 ( .IN1(n5769), .IN2(n4355), .S(n4326), .Q(n3649) );
  AO222X1 U3520 ( .IN1(N442), .IN2(n4322), .IN3(N378), .IN4(n4323), .IN5(n4324), .IN6(n4356), .Q(n3648) );
  MUX21X1 U3521 ( .IN1(n5770), .IN2(n4356), .S(n4326), .Q(n3647) );
  AO222X1 U3522 ( .IN1(N441), .IN2(n4322), .IN3(N377), .IN4(n4323), .IN5(n4324), .IN6(n4357), .Q(n3646) );
  MUX21X1 U3523 ( .IN1(n5771), .IN2(n4357), .S(n4326), .Q(n3645) );
  MUX21X1 U3524 ( .IN1(n5705), .IN2(ID_imm_offset[6]), .S(n4358), .Q(n3644) );
  AO22X1 U3525 ( .IN1(n4359), .IN2(n4253), .IN3(instruction[5]), .IN4(n4254), 
        .Q(n3643) );
  MUX21X1 U3526 ( .IN1(n4359), .IN2(ID_imm_offset[5]), .S(n4358), .Q(n3642) );
  AND2X1 U3527 ( .IN1(n4360), .IN2(n4261), .Q(n4358) );
  NAND4X0 U3528 ( .IN1(n4361), .IN2(n4362), .IN3(n4363), .IN4(n4364), .QN(
        n4261) );
  NAND2X0 U3529 ( .IN1(n4365), .IN2(n5736), .QN(n4363) );
  INVX0 U3530 ( .INP(N695), .ZN(n5736) );
  NAND2X0 U3531 ( .IN1(n4302), .IN2(n5739), .QN(n4362) );
  MUX21X1 U3532 ( .IN1(n4366), .IN2(n4367), .S(n3797), .Q(n4361) );
  NAND2X0 U3533 ( .IN1(n4252), .IN2(n4250), .QN(n4366) );
  NAND4X0 U3534 ( .IN1(n4368), .IN2(n3132), .IN3(n4250), .IN4(n4369), .QN(
        n4360) );
  INVX0 U3535 ( .INP(n5732), .ZN(n4359) );
  AO22X1 U3536 ( .IN1(n4370), .IN2(n4253), .IN3(instruction[4]), .IN4(n4254), 
        .Q(n3641) );
  MUX21X1 U3537 ( .IN1(n4371), .IN2(n4372), .S(N777), .Q(n3640) );
  AO22X1 U3538 ( .IN1(n4373), .IN2(n4370), .IN3(n4374), .IN4(n4243), .Q(n4372)
         );
  INVX0 U3539 ( .INP(n5733), .ZN(n4370) );
  AO22X1 U3540 ( .IN1(n5718), .IN2(n4253), .IN3(instruction[3]), .IN4(n4254), 
        .Q(n3639) );
  MUX21X1 U3541 ( .IN1(n4375), .IN2(n4376), .S(N777), .Q(n3638) );
  AO22X1 U3542 ( .IN1(n5718), .IN2(n4373), .IN3(n4374), .IN4(n4241), .Q(n4376)
         );
  AO22X1 U3543 ( .IN1(n4377), .IN2(n4253), .IN3(instruction[2]), .IN4(n4254), 
        .Q(n3637) );
  AO222X1 U3544 ( .IN1(n4378), .IN2(n4377), .IN3(n4379), .IN4(n5719), .IN5(
        n4380), .IN6(n4381), .Q(n3636) );
  AO222X1 U3545 ( .IN1(n4322), .IN2(n4243), .IN3(n4323), .IN4(n4377), .IN5(
        n4324), .IN6(n3880), .Q(n3635) );
  INVX0 U3546 ( .INP(n5729), .ZN(n4377) );
  MUX21X1 U3547 ( .IN1(n3808), .IN2(n3880), .S(n4254), .Q(n3634) );
  AO22X1 U3548 ( .IN1(n4382), .IN2(n4253), .IN3(instruction[1]), .IN4(n4254), 
        .Q(n3633) );
  AO222X1 U3549 ( .IN1(n4378), .IN2(n4382), .IN3(n4379), .IN4(n4260), .IN5(
        n4380), .IN6(n4383), .Q(n3632) );
  AO222X1 U3550 ( .IN1(n4322), .IN2(n4241), .IN3(n4323), .IN4(n4382), .IN5(
        n4324), .IN6(n3881), .Q(n3631) );
  INVX0 U3551 ( .INP(n5730), .ZN(n4382) );
  MUX21X1 U3552 ( .IN1(n3806), .IN2(n3881), .S(n4254), .Q(n3630) );
  AO22X1 U3553 ( .IN1(n5715), .IN2(n4253), .IN3(instruction[0]), .IN4(n4254), 
        .Q(n3629) );
  INVX0 U3554 ( .INP(reset_n), .ZN(n4253) );
  AO222X1 U3555 ( .IN1(n5715), .IN2(n4378), .IN3(n4379), .IN4(n5705), .IN5(
        n4380), .IN6(n4384), .Q(n3628) );
  AND2X1 U3556 ( .IN1(N773), .IN2(n4374), .Q(n4379) );
  AO21X1 U3557 ( .IN1(n4312), .IN2(n3131), .IN3(n4256), .Q(n4374) );
  NOR2X0 U3558 ( .IN1(n4364), .IN2(n4250), .QN(n4256) );
  NOR2X0 U3559 ( .IN1(n4380), .IN2(n4314), .QN(n4378) );
  INVX0 U3560 ( .INP(n4373), .ZN(n4314) );
  OA21X1 U3561 ( .IN1(n4367), .IN2(n4250), .IN3(n4364), .Q(n4373) );
  INVX0 U3562 ( .INP(n3131), .ZN(n4250) );
  INVX0 U3563 ( .INP(N773), .ZN(n4380) );
  AO222X1 U3564 ( .IN1(n4322), .IN2(n5719), .IN3(n5715), .IN4(n4323), .IN5(
        n4324), .IN6(n3809), .Q(n3627) );
  AOI21X1 U3565 ( .IN1(n4385), .IN2(n4364), .IN3(n4324), .QN(n4323) );
  INVX0 U3566 ( .INP(n4386), .ZN(n4324) );
  NAND2X0 U3567 ( .IN1(n4252), .IN2(n4248), .QN(n4364) );
  INVX0 U3568 ( .INP(n3130), .ZN(n4252) );
  MUX21X1 U3569 ( .IN1(n4320), .IN2(n4305), .S(n3132), .Q(n4385) );
  AND2X1 U3570 ( .IN1(n4387), .IN2(n4386), .Q(n4322) );
  AO221X1 U3571 ( .IN1(n4388), .IN2(n3131), .IN3(n4302), .IN4(n4389), .IN5(
        n4390), .Q(n4386) );
  MUX21X1 U3572 ( .IN1(n4312), .IN2(n4391), .S(n3797), .Q(n4390) );
  NOR2X0 U3573 ( .IN1(n3130), .IN2(n4365), .QN(n4391) );
  NOR2X0 U3574 ( .IN1(n3132), .IN2(n3131), .QN(n4365) );
  INVX0 U3575 ( .INP(n4367), .ZN(n4312) );
  NAND2X0 U3576 ( .IN1(n3132), .IN2(n3130), .QN(n4367) );
  NAND2X0 U3577 ( .IN1(n4248), .IN2(n5739), .QN(n4388) );
  INVX0 U3578 ( .INP(n3132), .ZN(n4248) );
  MUX21X1 U3579 ( .IN1(n3132), .IN2(n4392), .S(n4302), .Q(n4387) );
  INVX0 U3580 ( .INP(n4305), .ZN(n4302) );
  NAND2X0 U3581 ( .IN1(n3130), .IN2(n3131), .QN(n4305) );
  NOR2X0 U3582 ( .IN1(n3132), .IN2(n5739), .QN(n4392) );
  MUX21X1 U3583 ( .IN1(n3883), .IN2(n3809), .S(n4254), .Q(n3626) );
  NAND2X0 U3584 ( .IN1(n4393), .IN2(n4251), .QN(n3625) );
  MUX21X1 U3585 ( .IN1(n5709), .IN2(n5721), .S(reset_n), .Q(n4393) );
  NAND2X0 U3586 ( .IN1(n4394), .IN2(n4251), .QN(n3624) );
  MUX21X1 U3587 ( .IN1(n5707), .IN2(n5723), .S(reset_n), .Q(n4394) );
  NAND2X0 U3588 ( .IN1(n4395), .IN2(n4251), .QN(n3623) );
  MUX21X1 U3589 ( .IN1(n5708), .IN2(n5724), .S(reset_n), .Q(n4395) );
  NAND2X0 U3590 ( .IN1(n4396), .IN2(n4251), .QN(n3622) );
  NAND2X0 U3591 ( .IN1(reset_n), .IN2(n3842), .QN(n4251) );
  MUX21X1 U3592 ( .IN1(n5713), .IN2(\r150/A[3] ), .S(reset_n), .Q(n4396) );
  MUX21X1 U3593 ( .IN1(n3917), .IN2(n4397), .S(n4398), .Q(n3621) );
  NOR2X0 U3594 ( .IN1(n4399), .IN2(n4400), .QN(n4398) );
  AND3X1 U3595 ( .IN1(n4401), .IN2(n4402), .IN3(n4403), .Q(n4399) );
  MUX21X1 U3596 ( .IN1(n4404), .IN2(n4405), .S(n4406), .Q(n4403) );
  NAND2X0 U3597 ( .IN1(n4407), .IN2(n4408), .QN(n4405) );
  NAND3X0 U3598 ( .IN1(n5723), .IN2(n4409), .IN3(n4410), .QN(n4402) );
  AO21X1 U3599 ( .IN1(n4411), .IN2(n4412), .IN3(n4413), .Q(n4397) );
  NOR4X0 U3600 ( .IN1(n4414), .IN2(n4415), .IN3(n3804), .IN4(n3803), .QN(n4413) );
  NAND3X0 U3601 ( .IN1(n4416), .IN2(n3844), .IN3(n5723), .QN(n4414) );
  NAND3X0 U3602 ( .IN1(n4417), .IN2(n4401), .IN3(n4418), .QN(n4412) );
  AOI221X1 U3603 ( .IN1(n4419), .IN2(n4420), .IN3(n4421), .IN4(n3805), .IN5(
        n4422), .QN(n4401) );
  INVX0 U3604 ( .INP(n4423), .ZN(n4422) );
  AO222X1 U3605 ( .IN1(n4424), .IN2(n4425), .IN3(n4426), .IN4(n4427), .IN5(
        n4410), .IN6(n4428), .Q(n4421) );
  NOR2X0 U3606 ( .IN1(\r150/A[3] ), .IN2(n3843), .QN(n4426) );
  NOR2X0 U3607 ( .IN1(n5720), .IN2(n3844), .QN(n4424) );
  NOR2X0 U3608 ( .IN1(n3804), .IN2(n4429), .QN(n4419) );
  MUX21X1 U3609 ( .IN1(n4430), .IN2(n3847), .S(n4431), .Q(n4411) );
  MUX21X1 U3610 ( .IN1(n3879), .IN2(n314), .S(n4432), .Q(n3620) );
  MUX21X1 U3611 ( .IN1(n3878), .IN2(n313), .S(n4432), .Q(n3619) );
  MUX21X1 U3612 ( .IN1(n3877), .IN2(n312), .S(n4432), .Q(n3618) );
  MUX21X1 U3613 ( .IN1(n3876), .IN2(n311), .S(n4432), .Q(n3617) );
  MUX21X1 U3614 ( .IN1(n3875), .IN2(n310), .S(n4432), .Q(n3616) );
  MUX21X1 U3615 ( .IN1(n3874), .IN2(n309), .S(n4432), .Q(n3615) );
  MUX21X1 U3616 ( .IN1(n3873), .IN2(n308), .S(n4432), .Q(n3614) );
  MUX21X1 U3617 ( .IN1(n3872), .IN2(n307), .S(n4432), .Q(n3613) );
  MUX21X1 U3618 ( .IN1(n3871), .IN2(n306), .S(n4432), .Q(n3612) );
  MUX21X1 U3619 ( .IN1(n3870), .IN2(n305), .S(n4432), .Q(n3611) );
  MUX21X1 U3620 ( .IN1(n3869), .IN2(n304), .S(n4432), .Q(n3610) );
  MUX21X1 U3621 ( .IN1(n3868), .IN2(n303), .S(n4432), .Q(n3609) );
  MUX21X1 U3622 ( .IN1(n3867), .IN2(n302), .S(n4432), .Q(n3608) );
  MUX21X1 U3623 ( .IN1(n3866), .IN2(n301), .S(n4432), .Q(n3607) );
  MUX21X1 U3624 ( .IN1(n3865), .IN2(n300), .S(n4432), .Q(n3606) );
  MUX21X1 U3625 ( .IN1(n3864), .IN2(n299), .S(n4432), .Q(n3605) );
  MUX21X1 U3626 ( .IN1(n3863), .IN2(n298), .S(n4432), .Q(n3604) );
  MUX21X1 U3627 ( .IN1(n3862), .IN2(n297), .S(n4432), .Q(n3603) );
  MUX21X1 U3628 ( .IN1(n3861), .IN2(n296), .S(n4432), .Q(n3602) );
  MUX21X1 U3629 ( .IN1(n3860), .IN2(n295), .S(n4432), .Q(n3601) );
  MUX21X1 U3630 ( .IN1(n3859), .IN2(n294), .S(n4432), .Q(n3600) );
  MUX21X1 U3631 ( .IN1(n3858), .IN2(n293), .S(n4432), .Q(n3599) );
  MUX21X1 U3632 ( .IN1(n3857), .IN2(n292), .S(n4432), .Q(n3598) );
  MUX21X1 U3633 ( .IN1(n3856), .IN2(n291), .S(n4432), .Q(n3597) );
  MUX21X1 U3634 ( .IN1(n3855), .IN2(n290), .S(n4432), .Q(n3596) );
  MUX21X1 U3635 ( .IN1(n3854), .IN2(n289), .S(n4432), .Q(n3595) );
  MUX21X1 U3636 ( .IN1(n3853), .IN2(n288), .S(n4432), .Q(n3594) );
  MUX21X1 U3637 ( .IN1(n3852), .IN2(n287), .S(n4432), .Q(n3593) );
  MUX21X1 U3638 ( .IN1(n3851), .IN2(n286), .S(n4432), .Q(n3592) );
  MUX21X1 U3639 ( .IN1(n3850), .IN2(n285), .S(n4432), .Q(n3591) );
  MUX21X1 U3640 ( .IN1(n3849), .IN2(n284), .S(n4432), .Q(n3590) );
  MUX21X1 U3641 ( .IN1(n3848), .IN2(n283), .S(n4432), .Q(n3589) );
  AND2X1 U3642 ( .IN1(n3792), .IN2(reset_n), .Q(n4432) );
  NOR4X0 U3643 ( .IN1(n3842), .IN2(n4433), .IN3(n5722), .IN4(\r150/A[3] ), 
        .QN(n3792) );
  MUX21X1 U3644 ( .IN1(IF_PC[31]), .IN2(N344), .S(reset_n), .Q(n3588) );
  MUX21X1 U3645 ( .IN1(IF_PC[0]), .IN2(N313), .S(reset_n), .Q(n3587) );
  MUX21X1 U3646 ( .IN1(IF_PC[1]), .IN2(N314), .S(reset_n), .Q(n3586) );
  MUX21X1 U3647 ( .IN1(IF_PC[2]), .IN2(N315), .S(reset_n), .Q(n3585) );
  MUX21X1 U3648 ( .IN1(IF_PC[3]), .IN2(N316), .S(reset_n), .Q(n3584) );
  MUX21X1 U3649 ( .IN1(IF_PC[4]), .IN2(N317), .S(reset_n), .Q(n3583) );
  MUX21X1 U3650 ( .IN1(IF_PC[5]), .IN2(N318), .S(reset_n), .Q(n3582) );
  MUX21X1 U3651 ( .IN1(IF_PC[6]), .IN2(N319), .S(reset_n), .Q(n3581) );
  MUX21X1 U3652 ( .IN1(IF_PC[7]), .IN2(N320), .S(reset_n), .Q(n3580) );
  MUX21X1 U3653 ( .IN1(IF_PC[8]), .IN2(N321), .S(reset_n), .Q(n3579) );
  MUX21X1 U3654 ( .IN1(IF_PC[9]), .IN2(N322), .S(reset_n), .Q(n3578) );
  MUX21X1 U3655 ( .IN1(IF_PC[10]), .IN2(N323), .S(reset_n), .Q(n3577) );
  MUX21X1 U3656 ( .IN1(IF_PC[11]), .IN2(N324), .S(reset_n), .Q(n3576) );
  MUX21X1 U3657 ( .IN1(IF_PC[12]), .IN2(N325), .S(reset_n), .Q(n3575) );
  MUX21X1 U3658 ( .IN1(IF_PC[13]), .IN2(N326), .S(reset_n), .Q(n3574) );
  MUX21X1 U3659 ( .IN1(IF_PC[14]), .IN2(N327), .S(reset_n), .Q(n3573) );
  MUX21X1 U3660 ( .IN1(IF_PC[15]), .IN2(N328), .S(reset_n), .Q(n3572) );
  MUX21X1 U3661 ( .IN1(IF_PC[16]), .IN2(N329), .S(reset_n), .Q(n3571) );
  MUX21X1 U3662 ( .IN1(IF_PC[17]), .IN2(N330), .S(reset_n), .Q(n3570) );
  MUX21X1 U3663 ( .IN1(IF_PC[18]), .IN2(N331), .S(reset_n), .Q(n3569) );
  MUX21X1 U3664 ( .IN1(IF_PC[19]), .IN2(N332), .S(reset_n), .Q(n3568) );
  MUX21X1 U3665 ( .IN1(IF_PC[20]), .IN2(N333), .S(reset_n), .Q(n3567) );
  MUX21X1 U3666 ( .IN1(IF_PC[21]), .IN2(N334), .S(reset_n), .Q(n3566) );
  MUX21X1 U3667 ( .IN1(IF_PC[22]), .IN2(N335), .S(reset_n), .Q(n3565) );
  MUX21X1 U3668 ( .IN1(IF_PC[23]), .IN2(N336), .S(reset_n), .Q(n3564) );
  MUX21X1 U3669 ( .IN1(IF_PC[24]), .IN2(N337), .S(reset_n), .Q(n3563) );
  MUX21X1 U3670 ( .IN1(IF_PC[25]), .IN2(N338), .S(reset_n), .Q(n3562) );
  MUX21X1 U3671 ( .IN1(IF_PC[26]), .IN2(N339), .S(reset_n), .Q(n3561) );
  MUX21X1 U3672 ( .IN1(IF_PC[27]), .IN2(N340), .S(reset_n), .Q(n3560) );
  MUX21X1 U3673 ( .IN1(IF_PC[28]), .IN2(N341), .S(reset_n), .Q(n3559) );
  MUX21X1 U3674 ( .IN1(IF_PC[29]), .IN2(N342), .S(reset_n), .Q(n3558) );
  MUX21X1 U3675 ( .IN1(IF_PC[30]), .IN2(N343), .S(reset_n), .Q(n3557) );
  AO222X1 U3676 ( .IN1(n4434), .IN2(n283), .IN3(n4435), .IN4(N1244), .IN5(
        n4436), .IN6(SP[31]), .Q(n3556) );
  MUX21X1 U3677 ( .IN1(n3810), .IN2(n4437), .S(n4438), .Q(n3555) );
  MUX21X1 U3678 ( .IN1(data_address[0]), .IN2(n4437), .S(n4439), .Q(n3554) );
  AO222X1 U3679 ( .IN1(n4434), .IN2(n314), .IN3(N1213), .IN4(n4435), .IN5(
        n4436), .IN6(SP[0]), .Q(n3553) );
  AO222X1 U3680 ( .IN1(n4440), .IN2(n3810), .IN3(n4441), .IN4(n4437), .IN5(
        n4442), .IN6(n3916), .Q(n3552) );
  OR4X1 U3681 ( .IN1(n4443), .IN2(n4444), .IN3(n4445), .IN4(n4446), .Q(n4437)
         );
  AO221X1 U3682 ( .IN1(n4447), .IN2(n4448), .IN3(n4449), .IN4(n4450), .IN5(
        n4451), .Q(n4446) );
  AO22X1 U3683 ( .IN1(n4452), .IN2(n4453), .IN3(n4454), .IN4(n4455), .Q(n4451)
         );
  AO221X1 U3684 ( .IN1(n4456), .IN2(n4384), .IN3(n314), .IN4(n4457), .IN5(
        n4458), .Q(n4445) );
  AO222X1 U3685 ( .IN1(n4459), .IN2(n4460), .IN3(n4461), .IN4(n4462), .IN5(
        n4463), .IN6(n4464), .Q(n4458) );
  NOR2X0 U3686 ( .IN1(n3094), .IN2(n3062), .QN(n4461) );
  AO221X1 U3687 ( .IN1(N3556), .IN2(n4465), .IN3(N3827), .IN4(n4466), .IN5(
        n4467), .Q(n4444) );
  AO21X1 U3688 ( .IN1(N3688), .IN2(n4468), .IN3(n4469), .Q(n4467) );
  AO221X1 U3689 ( .IN1(N1148), .IN2(n4470), .IN3(N1213), .IN4(n4471), .IN5(
        n4472), .Q(n4443) );
  AO22X1 U3690 ( .IN1(N3724), .IN2(n4473), .IN3(N3791), .IN4(n4474), .Q(n4472)
         );
  MUX21X1 U3691 ( .IN1(n3811), .IN2(n4475), .S(n4438), .Q(n3551) );
  MUX21X1 U3692 ( .IN1(data_address[1]), .IN2(n4475), .S(n4439), .Q(n3550) );
  AO222X1 U3693 ( .IN1(n4434), .IN2(n313), .IN3(N1214), .IN4(n4435), .IN5(
        n4436), .IN6(SP[1]), .Q(n3549) );
  AO222X1 U3694 ( .IN1(n4440), .IN2(n3811), .IN3(n4441), .IN4(n4475), .IN5(
        n4442), .IN6(n3915), .Q(n3548) );
  OR4X1 U3695 ( .IN1(n4476), .IN2(n4477), .IN3(n4478), .IN4(n4479), .Q(n4475)
         );
  AO221X1 U3696 ( .IN1(n4447), .IN2(n4453), .IN3(n4452), .IN4(n4455), .IN5(
        n4480), .Q(n4479) );
  AO22X1 U3697 ( .IN1(n313), .IN2(n4457), .IN3(n4456), .IN4(n4383), .Q(n4480)
         );
  AO221X1 U3698 ( .IN1(n4454), .IN2(n4464), .IN3(n4463), .IN4(n4481), .IN5(
        n4482), .Q(n4478) );
  AO222X1 U3699 ( .IN1(n4449), .IN2(n4460), .IN3(n4483), .IN4(n4462), .IN5(
        n4459), .IN6(n4484), .Q(n4482) );
  NOR2X0 U3700 ( .IN1(n3093), .IN2(n3060), .QN(n4483) );
  AO222X1 U3701 ( .IN1(n4485), .IN2(n4486), .IN3(n4487), .IN4(n4488), .IN5(
        n4489), .IN6(n4490), .Q(n4460) );
  AO221X1 U3702 ( .IN1(N3557), .IN2(n4465), .IN3(N3828), .IN4(n4466), .IN5(
        n4491), .Q(n4477) );
  AO21X1 U3703 ( .IN1(N3689), .IN2(n4468), .IN3(n4469), .Q(n4491) );
  AO221X1 U3704 ( .IN1(N1149), .IN2(n4470), .IN3(N1214), .IN4(n4471), .IN5(
        n4492), .Q(n4476) );
  AO22X1 U3705 ( .IN1(N3725), .IN2(n4473), .IN3(N3792), .IN4(n4474), .Q(n4492)
         );
  MUX21X1 U3706 ( .IN1(n3812), .IN2(n4493), .S(n4438), .Q(n3547) );
  MUX21X1 U3707 ( .IN1(data_address[2]), .IN2(n4493), .S(n4439), .Q(n3546) );
  AO222X1 U3708 ( .IN1(n4434), .IN2(n312), .IN3(N1215), .IN4(n4435), .IN5(
        n4436), .IN6(SP[2]), .Q(n3545) );
  AO222X1 U3709 ( .IN1(n4440), .IN2(n3812), .IN3(n4441), .IN4(n4493), .IN5(
        n4442), .IN6(n3914), .Q(n3544) );
  OR4X1 U3710 ( .IN1(n4494), .IN2(n4495), .IN3(n4496), .IN4(n4497), .Q(n4493)
         );
  AO221X1 U3711 ( .IN1(n312), .IN2(n4457), .IN3(n4447), .IN4(n4455), .IN5(
        n4498), .Q(n4497) );
  AO22X1 U3712 ( .IN1(n4456), .IN2(n4381), .IN3(n4463), .IN4(n4499), .Q(n4498)
         );
  AO221X1 U3713 ( .IN1(n4452), .IN2(n4464), .IN3(n4454), .IN4(n4481), .IN5(
        n4500), .Q(n4496) );
  AO222X1 U3714 ( .IN1(n4449), .IN2(n4484), .IN3(n4501), .IN4(n4462), .IN5(
        n4459), .IN6(n4487), .Q(n4500) );
  NOR2X0 U3715 ( .IN1(n3092), .IN2(n3058), .QN(n4501) );
  AO222X1 U3716 ( .IN1(n4502), .IN2(n4488), .IN3(n4485), .IN4(n4487), .IN5(
        n4489), .IN6(n4486), .Q(n4484) );
  AO221X1 U3717 ( .IN1(N3558), .IN2(n4465), .IN3(N3829), .IN4(n4466), .IN5(
        n4503), .Q(n4495) );
  AO21X1 U3718 ( .IN1(N3690), .IN2(n4468), .IN3(n4469), .Q(n4503) );
  AO221X1 U3719 ( .IN1(N3793), .IN2(n4474), .IN3(N3726), .IN4(n4473), .IN5(
        n4504), .Q(n4494) );
  AO222X1 U3720 ( .IN1(N1215), .IN2(n4471), .IN3(N1150), .IN4(n4470), .IN5(
        N1183), .IN6(n4505), .Q(n4504) );
  MUX21X1 U3721 ( .IN1(n3813), .IN2(n4506), .S(n4438), .Q(n3543) );
  MUX21X1 U3722 ( .IN1(data_address[3]), .IN2(n4506), .S(n4439), .Q(n3542) );
  AO222X1 U3723 ( .IN1(n4434), .IN2(n311), .IN3(N1216), .IN4(n4435), .IN5(
        n4436), .IN6(SP[3]), .Q(n3541) );
  AO222X1 U3724 ( .IN1(n4440), .IN2(n3813), .IN3(n4441), .IN4(n4506), .IN5(
        n4442), .IN6(n3913), .Q(n3540) );
  OR4X1 U3725 ( .IN1(n4507), .IN2(n4508), .IN3(n4509), .IN4(n4510), .Q(n4506)
         );
  AO221X1 U3726 ( .IN1(n4454), .IN2(n4499), .IN3(n4463), .IN4(n4511), .IN5(
        n4512), .Q(n4510) );
  AO22X1 U3727 ( .IN1(n311), .IN2(n4457), .IN3(n4456), .IN4(n4375), .Q(n4512)
         );
  AO221X1 U3728 ( .IN1(n4459), .IN2(n4502), .IN3(n4452), .IN4(n4481), .IN5(
        n4513), .Q(n4509) );
  AO222X1 U3729 ( .IN1(n4449), .IN2(n4487), .IN3(n4514), .IN4(n4462), .IN5(
        n4447), .IN6(n4464), .Q(n4513) );
  AO222X1 U3730 ( .IN1(n4515), .IN2(n4516), .IN3(n4499), .IN4(n4488), .IN5(
        n4517), .IN6(n4518), .Q(n4464) );
  NOR2X0 U3731 ( .IN1(n3091), .IN2(n3056), .QN(n4514) );
  AO222X1 U3732 ( .IN1(n4519), .IN2(n4520), .IN3(n4521), .IN4(n4522), .IN5(
        n4523), .IN6(n4524), .Q(n4487) );
  AO221X1 U3733 ( .IN1(N3559), .IN2(n4465), .IN3(N3830), .IN4(n4466), .IN5(
        n4525), .Q(n4508) );
  AO21X1 U3734 ( .IN1(N3691), .IN2(n4468), .IN3(n4469), .Q(n4525) );
  AO221X1 U3735 ( .IN1(N3794), .IN2(n4474), .IN3(N3727), .IN4(n4473), .IN5(
        n4526), .Q(n4507) );
  AO222X1 U3736 ( .IN1(N1216), .IN2(n4471), .IN3(N1151), .IN4(n4470), .IN5(
        N1184), .IN6(n4505), .Q(n4526) );
  MUX21X1 U3737 ( .IN1(n3814), .IN2(n4527), .S(n4438), .Q(n3539) );
  MUX21X1 U3738 ( .IN1(data_address[4]), .IN2(n4527), .S(n4439), .Q(n3538) );
  AO222X1 U3739 ( .IN1(n4434), .IN2(n310), .IN3(N1217), .IN4(n4435), .IN5(
        n4436), .IN6(SP[4]), .Q(n3537) );
  AO222X1 U3740 ( .IN1(n4440), .IN2(n3814), .IN3(n4441), .IN4(n4527), .IN5(
        n4442), .IN6(n3912), .Q(n3536) );
  OR4X1 U3741 ( .IN1(n4528), .IN2(n4529), .IN3(n4530), .IN4(n4531), .Q(n4527)
         );
  AO221X1 U3742 ( .IN1(n4454), .IN2(n4511), .IN3(n4456), .IN4(n4371), .IN5(
        n4532), .Q(n4531) );
  AO22X1 U3743 ( .IN1(n310), .IN2(n4457), .IN3(n4463), .IN4(n4533), .Q(n4532)
         );
  AO221X1 U3744 ( .IN1(n4447), .IN2(n4481), .IN3(n4452), .IN4(n4499), .IN5(
        n4534), .Q(n4530) );
  AO222X1 U3745 ( .IN1(n4459), .IN2(n4535), .IN3(n4536), .IN4(n4462), .IN5(
        n4449), .IN6(n4502), .Q(n4534) );
  AO222X1 U3746 ( .IN1(n4537), .IN2(n4522), .IN3(n4519), .IN4(n4521), .IN5(
        n4523), .IN6(n4520), .Q(n4502) );
  NOR2X0 U3747 ( .IN1(n3090), .IN2(n3054), .QN(n4536) );
  AO222X1 U3748 ( .IN1(n4511), .IN2(n4488), .IN3(n4517), .IN4(n4499), .IN5(
        n4515), .IN6(n4518), .Q(n4481) );
  AO221X1 U3749 ( .IN1(N3560), .IN2(n4465), .IN3(N3831), .IN4(n4466), .IN5(
        n4538), .Q(n4529) );
  AO21X1 U3750 ( .IN1(N3692), .IN2(n4468), .IN3(n4469), .Q(n4538) );
  AO221X1 U3751 ( .IN1(N3795), .IN2(n4474), .IN3(N3728), .IN4(n4473), .IN5(
        n4539), .Q(n4528) );
  AO222X1 U3752 ( .IN1(N1217), .IN2(n4471), .IN3(N1152), .IN4(n4470), .IN5(
        N1185), .IN6(n4505), .Q(n4539) );
  MUX21X1 U3753 ( .IN1(n3815), .IN2(n4540), .S(n4438), .Q(n3535) );
  MUX21X1 U3754 ( .IN1(data_address[5]), .IN2(n4540), .S(n4439), .Q(n3534) );
  AO222X1 U3755 ( .IN1(n4434), .IN2(n309), .IN3(N1218), .IN4(n4435), .IN5(
        n4436), .IN6(SP[5]), .Q(n3533) );
  AO222X1 U3756 ( .IN1(n4440), .IN2(n3815), .IN3(n4441), .IN4(n4540), .IN5(
        n4442), .IN6(n3911), .Q(n3532) );
  OR4X1 U3757 ( .IN1(n4541), .IN2(n4542), .IN3(n4543), .IN4(n4544), .Q(n4540)
         );
  AO221X1 U3758 ( .IN1(n4463), .IN2(n4545), .IN3(n309), .IN4(n4457), .IN5(
        n4546), .Q(n4544) );
  AO22X1 U3759 ( .IN1(n4454), .IN2(n4533), .IN3(n4456), .IN4(ID_imm_offset[5]), 
        .Q(n4546) );
  AO221X1 U3760 ( .IN1(n4459), .IN2(n4537), .IN3(n4452), .IN4(n4511), .IN5(
        n4547), .Q(n4543) );
  AO222X1 U3761 ( .IN1(n4449), .IN2(n4535), .IN3(n4548), .IN4(n4462), .IN5(
        n4447), .IN6(n4499), .Q(n4547) );
  AO222X1 U3762 ( .IN1(n4549), .IN2(n4550), .IN3(n4533), .IN4(n4522), .IN5(
        n4551), .IN6(n4552), .Q(n4499) );
  NOR2X0 U3763 ( .IN1(n3089), .IN2(n3052), .QN(n4548) );
  AO222X1 U3764 ( .IN1(n4519), .IN2(n4537), .IN3(n4523), .IN4(n4521), .IN5(
        n4553), .IN6(n4522), .Q(n4535) );
  AO222X1 U3765 ( .IN1(n4554), .IN2(n4555), .IN3(n4553), .IN4(n4556), .IN5(
        n4557), .IN6(n4558), .Q(n4521) );
  AO221X1 U3766 ( .IN1(N3561), .IN2(n4465), .IN3(N3832), .IN4(n4466), .IN5(
        n4559), .Q(n4542) );
  AO21X1 U3767 ( .IN1(N3693), .IN2(n4468), .IN3(n4469), .Q(n4559) );
  AO221X1 U3768 ( .IN1(N3796), .IN2(n4474), .IN3(N3729), .IN4(n4473), .IN5(
        n4560), .Q(n4541) );
  AO222X1 U3769 ( .IN1(N1218), .IN2(n4471), .IN3(N1153), .IN4(n4470), .IN5(
        N1186), .IN6(n4505), .Q(n4560) );
  MUX21X1 U3770 ( .IN1(n3816), .IN2(n4561), .S(n4438), .Q(n3531) );
  MUX21X1 U3771 ( .IN1(data_address[6]), .IN2(n4561), .S(n4439), .Q(n3530) );
  AO222X1 U3772 ( .IN1(n4434), .IN2(n308), .IN3(N1219), .IN4(n4435), .IN5(
        n4436), .IN6(SP[6]), .Q(n3529) );
  AO222X1 U3773 ( .IN1(n4440), .IN2(n3816), .IN3(n4441), .IN4(n4561), .IN5(
        n4442), .IN6(n3910), .Q(n3528) );
  OR4X1 U3774 ( .IN1(n4562), .IN2(n4563), .IN3(n4564), .IN4(n4565), .Q(n4561)
         );
  AO221X1 U3775 ( .IN1(n4452), .IN2(n4533), .IN3(n4454), .IN4(n4545), .IN5(
        n4566), .Q(n4565) );
  AO22X1 U3776 ( .IN1(n308), .IN2(n4457), .IN3(n4463), .IN4(n4567), .Q(n4566)
         );
  AO221X1 U3777 ( .IN1(n4459), .IN2(n4553), .IN3(n4456), .IN4(ID_imm_offset[6]), .IN5(n4568), .Q(n4564) );
  AO222X1 U3778 ( .IN1(n4449), .IN2(n4537), .IN3(n4569), .IN4(n4462), .IN5(
        n4447), .IN6(n4511), .Q(n4568) );
  AO222X1 U3779 ( .IN1(n4545), .IN2(n4522), .IN3(n4551), .IN4(n4533), .IN5(
        n4549), .IN6(n4552), .Q(n4511) );
  NOR2X0 U3780 ( .IN1(n3088), .IN2(n3050), .QN(n4569) );
  AO222X1 U3781 ( .IN1(n4570), .IN2(n4556), .IN3(n4554), .IN4(n4553), .IN5(
        n4557), .IN6(n4555), .Q(n4537) );
  AO221X1 U3782 ( .IN1(N3562), .IN2(n4465), .IN3(N3833), .IN4(n4466), .IN5(
        n4571), .Q(n4563) );
  AO21X1 U3783 ( .IN1(N3694), .IN2(n4468), .IN3(n4469), .Q(n4571) );
  AO221X1 U3784 ( .IN1(N3797), .IN2(n4474), .IN3(N3730), .IN4(n4473), .IN5(
        n4572), .Q(n4562) );
  AO222X1 U3785 ( .IN1(N1219), .IN2(n4471), .IN3(N1154), .IN4(n4470), .IN5(
        N1187), .IN6(n4505), .Q(n4572) );
  MUX21X1 U3786 ( .IN1(n3817), .IN2(n4573), .S(n4438), .Q(n3527) );
  MUX21X1 U3787 ( .IN1(data_address[7]), .IN2(n4573), .S(n4439), .Q(n3526) );
  AO222X1 U3788 ( .IN1(n4434), .IN2(n307), .IN3(N1220), .IN4(n4435), .IN5(
        n4436), .IN6(SP[7]), .Q(n3525) );
  AO222X1 U3789 ( .IN1(n4440), .IN2(n3817), .IN3(n4441), .IN4(n4573), .IN5(
        n4442), .IN6(n3909), .Q(n3524) );
  OR4X1 U3790 ( .IN1(n4574), .IN2(n4575), .IN3(n4576), .IN4(n4577), .Q(n4573)
         );
  AO221X1 U3791 ( .IN1(n4452), .IN2(n4545), .IN3(n4454), .IN4(n4567), .IN5(
        n4578), .Q(n4577) );
  AO22X1 U3792 ( .IN1(n307), .IN2(n4457), .IN3(n4463), .IN4(n4579), .Q(n4578)
         );
  AO221X1 U3793 ( .IN1(n4447), .IN2(n4533), .IN3(n4459), .IN4(n4570), .IN5(
        n4580), .Q(n4576) );
  AO222X1 U3794 ( .IN1(n4449), .IN2(n4553), .IN3(n4581), .IN4(n4462), .IN5(
        n4456), .IN6(ID_imm_offset[7]), .Q(n4580) );
  NOR3X0 U3795 ( .IN1(n3804), .IN2(n5721), .IN3(n4582), .QN(n4456) );
  NOR2X0 U3796 ( .IN1(n3087), .IN2(n3048), .QN(n4581) );
  AO222X1 U3797 ( .IN1(n4583), .IN2(n4584), .IN3(n4585), .IN4(n4586), .IN5(
        n4587), .IN6(n4588), .Q(n4553) );
  AO222X1 U3798 ( .IN1(n4589), .IN2(n4590), .IN3(n4567), .IN4(n4591), .IN5(
        n4592), .IN6(n4593), .Q(n4533) );
  AO221X1 U3799 ( .IN1(N3563), .IN2(n4465), .IN3(N3834), .IN4(n4466), .IN5(
        n4594), .Q(n4575) );
  AO21X1 U3800 ( .IN1(N3695), .IN2(n4468), .IN3(n4469), .Q(n4594) );
  AO221X1 U3801 ( .IN1(N3798), .IN2(n4474), .IN3(N3731), .IN4(n4473), .IN5(
        n4595), .Q(n4574) );
  AO222X1 U3802 ( .IN1(N1220), .IN2(n4471), .IN3(N1155), .IN4(n4470), .IN5(
        N1188), .IN6(n4505), .Q(n4595) );
  MUX21X1 U3803 ( .IN1(n3818), .IN2(n4596), .S(n4438), .Q(n3523) );
  MUX21X1 U3804 ( .IN1(data_address[8]), .IN2(n4596), .S(n4439), .Q(n3522) );
  AO222X1 U3805 ( .IN1(n4434), .IN2(n306), .IN3(N1221), .IN4(n4435), .IN5(
        n4436), .IN6(SP[8]), .Q(n3521) );
  AO222X1 U3806 ( .IN1(n4440), .IN2(n3818), .IN3(n4441), .IN4(n4596), .IN5(
        n4442), .IN6(n3908), .Q(n3520) );
  OR4X1 U3807 ( .IN1(n4597), .IN2(n4598), .IN3(n4599), .IN4(n4600), .Q(n4596)
         );
  AO221X1 U3808 ( .IN1(n4454), .IN2(n4579), .IN3(n4463), .IN4(n4601), .IN5(
        n4602), .Q(n4600) );
  AO22X1 U3809 ( .IN1(N1156), .IN2(n4470), .IN3(n306), .IN4(n4457), .Q(n4602)
         );
  AO221X1 U3810 ( .IN1(n4459), .IN2(n4585), .IN3(n4452), .IN4(n4567), .IN5(
        n4603), .Q(n4599) );
  AO222X1 U3811 ( .IN1(n4449), .IN2(n4570), .IN3(n4604), .IN4(n4462), .IN5(
        n4447), .IN6(n4545), .Q(n4603) );
  AO222X1 U3812 ( .IN1(n4579), .IN2(n4591), .IN3(n4592), .IN4(n4567), .IN5(
        n4589), .IN6(n4593), .Q(n4545) );
  NOR2X0 U3813 ( .IN1(n3086), .IN2(n3046), .QN(n4604) );
  AO222X1 U3814 ( .IN1(n4605), .IN2(n4586), .IN3(n4583), .IN4(n4585), .IN5(
        n4584), .IN6(n4588), .Q(n4570) );
  AO221X1 U3815 ( .IN1(N3564), .IN2(n4465), .IN3(N3835), .IN4(n4466), .IN5(
        n4606), .Q(n4598) );
  AO21X1 U3816 ( .IN1(N3696), .IN2(n4468), .IN3(n4469), .Q(n4606) );
  AO221X1 U3817 ( .IN1(N3799), .IN2(n4474), .IN3(N3732), .IN4(n4473), .IN5(
        n4607), .Q(n4597) );
  AO22X1 U3818 ( .IN1(N1189), .IN2(n4505), .IN3(N1221), .IN4(n4471), .Q(n4607)
         );
  MUX21X1 U3819 ( .IN1(n3819), .IN2(n4608), .S(n4438), .Q(n3519) );
  MUX21X1 U3820 ( .IN1(data_address[9]), .IN2(n4608), .S(n4439), .Q(n3518) );
  AO222X1 U3821 ( .IN1(n4434), .IN2(n305), .IN3(N1222), .IN4(n4435), .IN5(
        n4436), .IN6(SP[9]), .Q(n3517) );
  AO222X1 U3822 ( .IN1(n4440), .IN2(n3819), .IN3(n4441), .IN4(n4608), .IN5(
        n4442), .IN6(n3907), .Q(n3516) );
  OR4X1 U3823 ( .IN1(n4609), .IN2(n4610), .IN3(n4611), .IN4(n4612), .Q(n4608)
         );
  AO221X1 U3824 ( .IN1(n4454), .IN2(n4601), .IN3(n4463), .IN4(n4613), .IN5(
        n4614), .Q(n4612) );
  AO22X1 U3825 ( .IN1(N1157), .IN2(n4470), .IN3(n305), .IN4(n4457), .Q(n4614)
         );
  AO221X1 U3826 ( .IN1(n4459), .IN2(n4605), .IN3(n4452), .IN4(n4579), .IN5(
        n4615), .Q(n4611) );
  AO222X1 U3827 ( .IN1(n4449), .IN2(n4585), .IN3(n4616), .IN4(n4462), .IN5(
        n4447), .IN6(n4567), .Q(n4615) );
  AO222X1 U3828 ( .IN1(n4557), .IN2(n4617), .IN3(n4601), .IN4(n4618), .IN5(
        n4619), .IN6(n4620), .Q(n4567) );
  NOR2X0 U3829 ( .IN1(n3085), .IN2(n3044), .QN(n4616) );
  AO222X1 U3830 ( .IN1(n4621), .IN2(n4622), .IN3(n4623), .IN4(n4591), .IN5(
        n4624), .IN6(n4625), .Q(n4585) );
  AO221X1 U3831 ( .IN1(N3565), .IN2(n4465), .IN3(N3836), .IN4(n4466), .IN5(
        n4626), .Q(n4610) );
  AO21X1 U3832 ( .IN1(N3697), .IN2(n4468), .IN3(n4469), .Q(n4626) );
  AO221X1 U3833 ( .IN1(N3800), .IN2(n4474), .IN3(N3733), .IN4(n4473), .IN5(
        n4627), .Q(n4609) );
  AO22X1 U3834 ( .IN1(N1190), .IN2(n4505), .IN3(N1222), .IN4(n4471), .Q(n4627)
         );
  MUX21X1 U3835 ( .IN1(n3820), .IN2(n4628), .S(n4438), .Q(n3515) );
  MUX21X1 U3836 ( .IN1(data_address[10]), .IN2(n4628), .S(n4439), .Q(n3514) );
  AO222X1 U3837 ( .IN1(n4434), .IN2(n304), .IN3(N1223), .IN4(n4435), .IN5(
        n4436), .IN6(SP[10]), .Q(n3513) );
  AO222X1 U3838 ( .IN1(n4440), .IN2(n3820), .IN3(n4441), .IN4(n4628), .IN5(
        n4442), .IN6(n3906), .Q(n3512) );
  OR4X1 U3839 ( .IN1(n4629), .IN2(n4630), .IN3(n4631), .IN4(n4632), .Q(n4628)
         );
  AO221X1 U3840 ( .IN1(n4454), .IN2(n4613), .IN3(n4463), .IN4(n4633), .IN5(
        n4634), .Q(n4632) );
  AO22X1 U3841 ( .IN1(N1158), .IN2(n4470), .IN3(n304), .IN4(n4457), .Q(n4634)
         );
  AO221X1 U3842 ( .IN1(n4459), .IN2(n4623), .IN3(n4452), .IN4(n4601), .IN5(
        n4635), .Q(n4631) );
  AO222X1 U3843 ( .IN1(n4449), .IN2(n4605), .IN3(n4636), .IN4(n4462), .IN5(
        n4447), .IN6(n4579), .Q(n4635) );
  AO222X1 U3844 ( .IN1(n4613), .IN2(n4618), .IN3(n4619), .IN4(n4601), .IN5(
        n4557), .IN6(n4620), .Q(n4579) );
  NOR2X0 U3845 ( .IN1(n3084), .IN2(n3042), .QN(n4636) );
  AO222X1 U3846 ( .IN1(n4637), .IN2(n4591), .IN3(n4621), .IN4(n4623), .IN5(
        n4624), .IN6(n4622), .Q(n4605) );
  AO221X1 U3847 ( .IN1(N3566), .IN2(n4465), .IN3(N3837), .IN4(n4466), .IN5(
        n4638), .Q(n4630) );
  AO21X1 U3848 ( .IN1(N3698), .IN2(n4468), .IN3(n4469), .Q(n4638) );
  AO221X1 U3849 ( .IN1(N3801), .IN2(n4474), .IN3(N3734), .IN4(n4473), .IN5(
        n4639), .Q(n4629) );
  AO22X1 U3850 ( .IN1(N1191), .IN2(n4505), .IN3(N1223), .IN4(n4471), .Q(n4639)
         );
  MUX21X1 U3851 ( .IN1(n3821), .IN2(n4640), .S(n4438), .Q(n3511) );
  MUX21X1 U3852 ( .IN1(data_address[11]), .IN2(n4640), .S(n4439), .Q(n3510) );
  AO222X1 U3853 ( .IN1(n4434), .IN2(n303), .IN3(N1224), .IN4(n4435), .IN5(
        n4436), .IN6(SP[11]), .Q(n3509) );
  AO222X1 U3854 ( .IN1(n4440), .IN2(n3821), .IN3(n4441), .IN4(n4640), .IN5(
        n4442), .IN6(n3905), .Q(n3508) );
  OR4X1 U3855 ( .IN1(n4641), .IN2(n4642), .IN3(n4643), .IN4(n4644), .Q(n4640)
         );
  AO221X1 U3856 ( .IN1(n4454), .IN2(n4633), .IN3(n4463), .IN4(n4645), .IN5(
        n4646), .Q(n4644) );
  AO22X1 U3857 ( .IN1(N1159), .IN2(n4470), .IN3(n303), .IN4(n4457), .Q(n4646)
         );
  AO221X1 U3858 ( .IN1(n4459), .IN2(n4637), .IN3(n4452), .IN4(n4613), .IN5(
        n4647), .Q(n4643) );
  AO222X1 U3859 ( .IN1(n4449), .IN2(n4623), .IN3(n4648), .IN4(n4462), .IN5(
        n4447), .IN6(n4601), .Q(n4647) );
  AO222X1 U3860 ( .IN1(n4649), .IN2(n4650), .IN3(n4633), .IN4(n4651), .IN5(
        n4652), .IN6(n4653), .Q(n4601) );
  NOR2X0 U3861 ( .IN1(n3083), .IN2(n3040), .QN(n4648) );
  AO222X1 U3862 ( .IN1(n4654), .IN2(n4655), .IN3(n4656), .IN4(n4657), .IN5(
        n4658), .IN6(n4659), .Q(n4623) );
  AO221X1 U3863 ( .IN1(N3567), .IN2(n4465), .IN3(N3838), .IN4(n4466), .IN5(
        n4660), .Q(n4642) );
  AO21X1 U3864 ( .IN1(N3699), .IN2(n4468), .IN3(n4469), .Q(n4660) );
  AO221X1 U3865 ( .IN1(N3802), .IN2(n4474), .IN3(N3735), .IN4(n4473), .IN5(
        n4661), .Q(n4641) );
  AO22X1 U3866 ( .IN1(N1192), .IN2(n4505), .IN3(N1224), .IN4(n4471), .Q(n4661)
         );
  MUX21X1 U3867 ( .IN1(n3822), .IN2(n4662), .S(n4438), .Q(n3507) );
  MUX21X1 U3868 ( .IN1(data_address[12]), .IN2(n4662), .S(n4439), .Q(n3506) );
  AO222X1 U3869 ( .IN1(n4434), .IN2(n302), .IN3(N1225), .IN4(n4435), .IN5(
        n4436), .IN6(SP[12]), .Q(n3505) );
  AO222X1 U3870 ( .IN1(n4440), .IN2(n3822), .IN3(n4441), .IN4(n4662), .IN5(
        n4442), .IN6(n3904), .Q(n3504) );
  OR4X1 U3871 ( .IN1(n4663), .IN2(n4664), .IN3(n4665), .IN4(n4666), .Q(n4662)
         );
  AO221X1 U3872 ( .IN1(n4454), .IN2(n4645), .IN3(n4463), .IN4(n4667), .IN5(
        n4668), .Q(n4666) );
  AO22X1 U3873 ( .IN1(N1160), .IN2(n4470), .IN3(n302), .IN4(n4457), .Q(n4668)
         );
  AO221X1 U3874 ( .IN1(n4459), .IN2(n4657), .IN3(n4452), .IN4(n4633), .IN5(
        n4669), .Q(n4665) );
  AO222X1 U3875 ( .IN1(n4449), .IN2(n4637), .IN3(n4670), .IN4(n4462), .IN5(
        n4447), .IN6(n4613), .Q(n4669) );
  AO222X1 U3876 ( .IN1(n4645), .IN2(n4651), .IN3(n4652), .IN4(n4633), .IN5(
        n4649), .IN6(n4653), .Q(n4613) );
  NOR2X0 U3877 ( .IN1(n3082), .IN2(n3038), .QN(n4670) );
  AO222X1 U3878 ( .IN1(n4656), .IN2(n4671), .IN3(n4654), .IN4(n4657), .IN5(
        n4658), .IN6(n4655), .Q(n4637) );
  AO221X1 U3879 ( .IN1(N3568), .IN2(n4465), .IN3(N3839), .IN4(n4466), .IN5(
        n4672), .Q(n4664) );
  AO21X1 U3880 ( .IN1(N3700), .IN2(n4468), .IN3(n4469), .Q(n4672) );
  AO221X1 U3881 ( .IN1(N3803), .IN2(n4474), .IN3(N3736), .IN4(n4473), .IN5(
        n4673), .Q(n4663) );
  AO22X1 U3882 ( .IN1(N1193), .IN2(n4505), .IN3(N1225), .IN4(n4471), .Q(n4673)
         );
  MUX21X1 U3883 ( .IN1(n3823), .IN2(n4674), .S(n4438), .Q(n3503) );
  MUX21X1 U3884 ( .IN1(data_address[13]), .IN2(n4674), .S(n4439), .Q(n3502) );
  AO222X1 U3885 ( .IN1(n4434), .IN2(n301), .IN3(N1226), .IN4(n4435), .IN5(
        n4436), .IN6(SP[13]), .Q(n3501) );
  AO222X1 U3886 ( .IN1(n4440), .IN2(n3823), .IN3(n4441), .IN4(n4674), .IN5(
        n4442), .IN6(n3903), .Q(n3500) );
  OR4X1 U3887 ( .IN1(n4675), .IN2(n4676), .IN3(n4677), .IN4(n4678), .Q(n4674)
         );
  AO221X1 U3888 ( .IN1(n4454), .IN2(n4667), .IN3(n4463), .IN4(n4679), .IN5(
        n4680), .Q(n4678) );
  AO22X1 U3889 ( .IN1(N1161), .IN2(n4470), .IN3(n301), .IN4(n4457), .Q(n4680)
         );
  AO221X1 U3890 ( .IN1(n4459), .IN2(n4671), .IN3(n4452), .IN4(n4645), .IN5(
        n4681), .Q(n4677) );
  AO222X1 U3891 ( .IN1(n4449), .IN2(n4657), .IN3(n4682), .IN4(n4462), .IN5(
        n4447), .IN6(n4633), .Q(n4681) );
  AO222X1 U3892 ( .IN1(n4683), .IN2(n4684), .IN3(n4667), .IN4(n4685), .IN5(
        n4686), .IN6(n4687), .Q(n4633) );
  NOR2X0 U3893 ( .IN1(n3081), .IN2(n3036), .QN(n4682) );
  AO222X1 U3894 ( .IN1(n4688), .IN2(n4689), .IN3(n4690), .IN4(n4691), .IN5(
        n4692), .IN6(n4693), .Q(n4657) );
  AO221X1 U3895 ( .IN1(N3569), .IN2(n4465), .IN3(N3840), .IN4(n4466), .IN5(
        n4694), .Q(n4676) );
  AO21X1 U3896 ( .IN1(N3701), .IN2(n4468), .IN3(n4469), .Q(n4694) );
  AO221X1 U3897 ( .IN1(N3804), .IN2(n4474), .IN3(N3737), .IN4(n4473), .IN5(
        n4695), .Q(n4675) );
  AO22X1 U3898 ( .IN1(N1194), .IN2(n4505), .IN3(N1226), .IN4(n4471), .Q(n4695)
         );
  MUX21X1 U3899 ( .IN1(n3824), .IN2(n4696), .S(n4438), .Q(n3499) );
  MUX21X1 U3900 ( .IN1(data_address[14]), .IN2(n4696), .S(n4439), .Q(n3498) );
  AO222X1 U3901 ( .IN1(n4434), .IN2(n300), .IN3(N1227), .IN4(n4435), .IN5(
        n4436), .IN6(SP[14]), .Q(n3497) );
  AO222X1 U3902 ( .IN1(n4440), .IN2(n3824), .IN3(n4441), .IN4(n4696), .IN5(
        n4442), .IN6(n3902), .Q(n3496) );
  OR4X1 U3903 ( .IN1(n4697), .IN2(n4698), .IN3(n4699), .IN4(n4700), .Q(n4696)
         );
  AO221X1 U3904 ( .IN1(n4454), .IN2(n4679), .IN3(n4463), .IN4(n4701), .IN5(
        n4702), .Q(n4700) );
  AO22X1 U3905 ( .IN1(N1162), .IN2(n4470), .IN3(n300), .IN4(n4457), .Q(n4702)
         );
  AO221X1 U3906 ( .IN1(n4459), .IN2(n4703), .IN3(n4452), .IN4(n4667), .IN5(
        n4704), .Q(n4699) );
  AO222X1 U3907 ( .IN1(n4449), .IN2(n4671), .IN3(n4705), .IN4(n4462), .IN5(
        n4447), .IN6(n4645), .Q(n4704) );
  AO222X1 U3908 ( .IN1(n4679), .IN2(n4685), .IN3(n4686), .IN4(n4667), .IN5(
        n4683), .IN6(n4687), .Q(n4645) );
  NOR2X0 U3909 ( .IN1(n3080), .IN2(n3034), .QN(n4705) );
  AO222X1 U3910 ( .IN1(n4706), .IN2(n4691), .IN3(n4688), .IN4(n4690), .IN5(
        n4692), .IN6(n4689), .Q(n4671) );
  AO221X1 U3911 ( .IN1(N3570), .IN2(n4465), .IN3(N3841), .IN4(n4466), .IN5(
        n4707), .Q(n4698) );
  AO21X1 U3912 ( .IN1(N3702), .IN2(n4468), .IN3(n4469), .Q(n4707) );
  AO221X1 U3913 ( .IN1(N3805), .IN2(n4474), .IN3(N3738), .IN4(n4473), .IN5(
        n4708), .Q(n4697) );
  AO22X1 U3914 ( .IN1(N1195), .IN2(n4505), .IN3(N1227), .IN4(n4471), .Q(n4708)
         );
  MUX21X1 U3915 ( .IN1(n3825), .IN2(n4709), .S(n4438), .Q(n3495) );
  MUX21X1 U3916 ( .IN1(data_address[15]), .IN2(n4709), .S(n4439), .Q(n3494) );
  AO222X1 U3917 ( .IN1(n4434), .IN2(n299), .IN3(N1228), .IN4(n4435), .IN5(
        n4436), .IN6(SP[15]), .Q(n3493) );
  AO222X1 U3918 ( .IN1(n4440), .IN2(n3825), .IN3(n4441), .IN4(n4709), .IN5(
        n4442), .IN6(n3901), .Q(n3492) );
  OR4X1 U3919 ( .IN1(n4710), .IN2(n4711), .IN3(n4712), .IN4(n4713), .Q(n4709)
         );
  AO221X1 U3920 ( .IN1(n4454), .IN2(n4701), .IN3(n4463), .IN4(n4714), .IN5(
        n4715), .Q(n4713) );
  AO22X1 U3921 ( .IN1(N1163), .IN2(n4470), .IN3(n299), .IN4(n4457), .Q(n4715)
         );
  AO221X1 U3922 ( .IN1(n4459), .IN2(n4706), .IN3(n4452), .IN4(n4679), .IN5(
        n4716), .Q(n4712) );
  AO222X1 U3923 ( .IN1(n4449), .IN2(n4703), .IN3(n4717), .IN4(n4462), .IN5(
        n4447), .IN6(n4667), .Q(n4716) );
  AO222X1 U3924 ( .IN1(n4718), .IN2(n4719), .IN3(n4701), .IN4(n4720), .IN5(
        n4721), .IN6(n4722), .Q(n4667) );
  NOR2X0 U3925 ( .IN1(n3079), .IN2(n3032), .QN(n4717) );
  AO222X1 U3926 ( .IN1(n4688), .IN2(n4706), .IN3(n4692), .IN4(n4690), .IN5(
        n4723), .IN6(n4691), .Q(n4703) );
  AO222X1 U3927 ( .IN1(n4724), .IN2(n4725), .IN3(n4723), .IN4(n4726), .IN5(
        n4727), .IN6(n4728), .Q(n4690) );
  AO221X1 U3928 ( .IN1(N3571), .IN2(n4465), .IN3(N3842), .IN4(n4466), .IN5(
        n4729), .Q(n4711) );
  AO21X1 U3929 ( .IN1(N3703), .IN2(n4468), .IN3(n4469), .Q(n4729) );
  AO221X1 U3930 ( .IN1(N3806), .IN2(n4474), .IN3(N3739), .IN4(n4473), .IN5(
        n4730), .Q(n4710) );
  AO22X1 U3931 ( .IN1(N1196), .IN2(n4505), .IN3(N1228), .IN4(n4471), .Q(n4730)
         );
  MUX21X1 U3932 ( .IN1(n3826), .IN2(n4731), .S(n4438), .Q(n3491) );
  MUX21X1 U3933 ( .IN1(data_address[16]), .IN2(n4731), .S(n4439), .Q(n3490) );
  AO222X1 U3934 ( .IN1(n4434), .IN2(n298), .IN3(N1229), .IN4(n4435), .IN5(
        n4436), .IN6(SP[16]), .Q(n3489) );
  AO222X1 U3935 ( .IN1(n4440), .IN2(n3826), .IN3(n4441), .IN4(n4731), .IN5(
        n4442), .IN6(n3900), .Q(n3488) );
  OR4X1 U3936 ( .IN1(n4732), .IN2(n4733), .IN3(n4734), .IN4(n4735), .Q(n4731)
         );
  AO221X1 U3937 ( .IN1(n4454), .IN2(n4714), .IN3(n4463), .IN4(n4736), .IN5(
        n4737), .Q(n4735) );
  AO22X1 U3938 ( .IN1(N1164), .IN2(n4470), .IN3(n298), .IN4(n4457), .Q(n4737)
         );
  AO221X1 U3939 ( .IN1(n4459), .IN2(n4723), .IN3(n4452), .IN4(n4701), .IN5(
        n4738), .Q(n4734) );
  AO222X1 U3940 ( .IN1(n4449), .IN2(n4706), .IN3(n4739), .IN4(n4462), .IN5(
        n4447), .IN6(n4679), .Q(n4738) );
  AO222X1 U3941 ( .IN1(n4714), .IN2(n4720), .IN3(n4721), .IN4(n4701), .IN5(
        n4718), .IN6(n4722), .Q(n4679) );
  NOR2X0 U3942 ( .IN1(n3078), .IN2(n3030), .QN(n4739) );
  AO222X1 U3943 ( .IN1(n4740), .IN2(n4726), .IN3(n4724), .IN4(n4723), .IN5(
        n4727), .IN6(n4725), .Q(n4706) );
  AO221X1 U3944 ( .IN1(N3572), .IN2(n4465), .IN3(N3843), .IN4(n4466), .IN5(
        n4741), .Q(n4733) );
  AO21X1 U3945 ( .IN1(N3704), .IN2(n4468), .IN3(n4469), .Q(n4741) );
  AO221X1 U3946 ( .IN1(N3807), .IN2(n4474), .IN3(N3740), .IN4(n4473), .IN5(
        n4742), .Q(n4732) );
  AO22X1 U3947 ( .IN1(N1197), .IN2(n4505), .IN3(N1229), .IN4(n4471), .Q(n4742)
         );
  MUX21X1 U3948 ( .IN1(n3827), .IN2(n4743), .S(n4438), .Q(n3487) );
  MUX21X1 U3949 ( .IN1(data_address[17]), .IN2(n4743), .S(n4439), .Q(n3486) );
  AO222X1 U3950 ( .IN1(n4434), .IN2(n297), .IN3(N1230), .IN4(n4435), .IN5(
        n4436), .IN6(SP[17]), .Q(n3485) );
  AO222X1 U3951 ( .IN1(n4440), .IN2(n3827), .IN3(n4441), .IN4(n4743), .IN5(
        n4442), .IN6(n3899), .Q(n3484) );
  OR4X1 U3952 ( .IN1(n4744), .IN2(n4745), .IN3(n4746), .IN4(n4747), .Q(n4743)
         );
  AO221X1 U3953 ( .IN1(n4454), .IN2(n4736), .IN3(n4463), .IN4(n4748), .IN5(
        n4749), .Q(n4747) );
  AO22X1 U3954 ( .IN1(N1165), .IN2(n4470), .IN3(n297), .IN4(n4457), .Q(n4749)
         );
  AO221X1 U3955 ( .IN1(n4459), .IN2(n4750), .IN3(n4452), .IN4(n4714), .IN5(
        n4751), .Q(n4746) );
  AO222X1 U3956 ( .IN1(n4449), .IN2(n4723), .IN3(n4752), .IN4(n4462), .IN5(
        n4447), .IN6(n4701), .Q(n4751) );
  AO222X1 U3957 ( .IN1(n4753), .IN2(n4754), .IN3(n4736), .IN4(n4755), .IN5(
        n4756), .IN6(n4757), .Q(n4701) );
  NOR2X0 U3958 ( .IN1(n3077), .IN2(n3028), .QN(n4752) );
  AO222X1 U3959 ( .IN1(n4758), .IN2(n4759), .IN3(n4760), .IN4(n4761), .IN5(
        n4762), .IN6(n4763), .Q(n4723) );
  AO221X1 U3960 ( .IN1(N3573), .IN2(n4465), .IN3(N3844), .IN4(n4466), .IN5(
        n4764), .Q(n4745) );
  AO21X1 U3961 ( .IN1(N3705), .IN2(n4468), .IN3(n4469), .Q(n4764) );
  AO221X1 U3962 ( .IN1(N3808), .IN2(n4474), .IN3(N3741), .IN4(n4473), .IN5(
        n4765), .Q(n4744) );
  AO22X1 U3963 ( .IN1(N1198), .IN2(n4505), .IN3(N1230), .IN4(n4471), .Q(n4765)
         );
  MUX21X1 U3964 ( .IN1(n3828), .IN2(n4766), .S(n4438), .Q(n3483) );
  MUX21X1 U3965 ( .IN1(data_address[18]), .IN2(n4766), .S(n4439), .Q(n3482) );
  AO222X1 U3966 ( .IN1(n4434), .IN2(n296), .IN3(N1231), .IN4(n4435), .IN5(
        n4436), .IN6(SP[18]), .Q(n3481) );
  AO222X1 U3967 ( .IN1(n4440), .IN2(n3828), .IN3(n4441), .IN4(n4766), .IN5(
        n4442), .IN6(n3898), .Q(n3480) );
  OR4X1 U3968 ( .IN1(n4767), .IN2(n4768), .IN3(n4769), .IN4(n4770), .Q(n4766)
         );
  AO221X1 U3969 ( .IN1(n4454), .IN2(n4748), .IN3(n4463), .IN4(n4771), .IN5(
        n4772), .Q(n4770) );
  AO22X1 U3970 ( .IN1(N1166), .IN2(n4470), .IN3(n296), .IN4(n4457), .Q(n4772)
         );
  AO221X1 U3971 ( .IN1(n4459), .IN2(n4773), .IN3(n4452), .IN4(n4736), .IN5(
        n4774), .Q(n4769) );
  AO222X1 U3972 ( .IN1(n4449), .IN2(n4750), .IN3(n4775), .IN4(n4462), .IN5(
        n4447), .IN6(n4714), .Q(n4774) );
  AO222X1 U3973 ( .IN1(n4748), .IN2(n4755), .IN3(n4756), .IN4(n4736), .IN5(
        n4753), .IN6(n4757), .Q(n4714) );
  NOR2X0 U3974 ( .IN1(n3076), .IN2(n3026), .QN(n4775) );
  AO21X1 U3975 ( .IN1(n4776), .IN2(n4691), .IN3(n4740), .Q(n4750) );
  AO222X1 U3976 ( .IN1(n4777), .IN2(n4761), .IN3(n4758), .IN4(n4760), .IN5(
        n4762), .IN6(n4759), .Q(n4740) );
  AO221X1 U3977 ( .IN1(N3574), .IN2(n4465), .IN3(N3845), .IN4(n4466), .IN5(
        n4778), .Q(n4768) );
  AO21X1 U3978 ( .IN1(N3706), .IN2(n4468), .IN3(n4469), .Q(n4778) );
  AO221X1 U3979 ( .IN1(N3809), .IN2(n4474), .IN3(N3742), .IN4(n4473), .IN5(
        n4779), .Q(n4767) );
  AO22X1 U3980 ( .IN1(N1199), .IN2(n4505), .IN3(N1231), .IN4(n4471), .Q(n4779)
         );
  MUX21X1 U3981 ( .IN1(n3829), .IN2(n4780), .S(n4438), .Q(n3479) );
  MUX21X1 U3982 ( .IN1(data_address[19]), .IN2(n4780), .S(n4439), .Q(n3478) );
  AO222X1 U3983 ( .IN1(n4434), .IN2(n295), .IN3(N1232), .IN4(n4435), .IN5(
        n4436), .IN6(SP[19]), .Q(n3477) );
  AO222X1 U3984 ( .IN1(n4440), .IN2(n3829), .IN3(n4441), .IN4(n4780), .IN5(
        n4442), .IN6(n3897), .Q(n3476) );
  OR4X1 U3985 ( .IN1(n4781), .IN2(n4782), .IN3(n4783), .IN4(n4784), .Q(n4780)
         );
  AO221X1 U3986 ( .IN1(n4454), .IN2(n4771), .IN3(n4463), .IN4(n4785), .IN5(
        n4786), .Q(n4784) );
  AO22X1 U3987 ( .IN1(N1167), .IN2(n4470), .IN3(n295), .IN4(n4457), .Q(n4786)
         );
  AO221X1 U3988 ( .IN1(n4459), .IN2(n4776), .IN3(n4452), .IN4(n4748), .IN5(
        n4787), .Q(n4783) );
  AO222X1 U3989 ( .IN1(n4449), .IN2(n4773), .IN3(n4788), .IN4(n4462), .IN5(
        n4447), .IN6(n4736), .Q(n4787) );
  AO222X1 U3990 ( .IN1(n4789), .IN2(n4790), .IN3(n4771), .IN4(n4791), .IN5(
        n4792), .IN6(n4793), .Q(n4736) );
  NOR2X0 U3991 ( .IN1(n3075), .IN2(n3024), .QN(n4788) );
  AO221X1 U3992 ( .IN1(n4794), .IN2(n4761), .IN3(n4795), .IN4(n4691), .IN5(
        n4796), .Q(n4773) );
  AO22X1 U3993 ( .IN1(n4758), .IN2(n4777), .IN3(n4762), .IN4(n4760), .Q(n4796)
         );
  AO222X1 U3994 ( .IN1(n4797), .IN2(n4798), .IN3(n4799), .IN4(n4720), .IN5(
        n4753), .IN6(n4800), .Q(n4760) );
  AO221X1 U3995 ( .IN1(N3575), .IN2(n4465), .IN3(N3846), .IN4(n4466), .IN5(
        n4801), .Q(n4782) );
  AO21X1 U3996 ( .IN1(N3707), .IN2(n4468), .IN3(n4469), .Q(n4801) );
  AO221X1 U3997 ( .IN1(N3810), .IN2(n4474), .IN3(N3743), .IN4(n4473), .IN5(
        n4802), .Q(n4781) );
  AO22X1 U3998 ( .IN1(N1200), .IN2(n4505), .IN3(N1232), .IN4(n4471), .Q(n4802)
         );
  MUX21X1 U3999 ( .IN1(n3830), .IN2(n4803), .S(n4438), .Q(n3475) );
  MUX21X1 U4000 ( .IN1(data_address[20]), .IN2(n4803), .S(n4439), .Q(n3474) );
  AO222X1 U4001 ( .IN1(n4434), .IN2(n294), .IN3(N1233), .IN4(n4435), .IN5(
        n4436), .IN6(SP[20]), .Q(n3473) );
  AO222X1 U4002 ( .IN1(n4440), .IN2(n3830), .IN3(n4441), .IN4(n4803), .IN5(
        n4442), .IN6(n3896), .Q(n3472) );
  OR4X1 U4003 ( .IN1(n4804), .IN2(n4805), .IN3(n4806), .IN4(n4807), .Q(n4803)
         );
  AO221X1 U4004 ( .IN1(n4454), .IN2(n4785), .IN3(n4463), .IN4(n4808), .IN5(
        n4809), .Q(n4807) );
  AO22X1 U4005 ( .IN1(N1168), .IN2(n4470), .IN3(n294), .IN4(n4457), .Q(n4809)
         );
  AO221X1 U4006 ( .IN1(n4459), .IN2(n4795), .IN3(n4452), .IN4(n4771), .IN5(
        n4810), .Q(n4806) );
  AO222X1 U4007 ( .IN1(n4449), .IN2(n4776), .IN3(n4811), .IN4(n4462), .IN5(
        n4447), .IN6(n4748), .Q(n4810) );
  AO222X1 U4008 ( .IN1(n4785), .IN2(n4791), .IN3(n4792), .IN4(n4771), .IN5(
        n4789), .IN6(n4793), .Q(n4748) );
  NOR2X0 U4009 ( .IN1(n3074), .IN2(n3022), .QN(n4811) );
  AO222X1 U4010 ( .IN1(n4758), .IN2(n4794), .IN3(n4762), .IN4(n4777), .IN5(
        n4812), .IN6(n4761), .Q(n4776) );
  AO222X1 U4011 ( .IN1(n4813), .IN2(n4720), .IN3(n4797), .IN4(n4799), .IN5(
        n4753), .IN6(n4798), .Q(n4777) );
  AO221X1 U4012 ( .IN1(N3576), .IN2(n4465), .IN3(N3847), .IN4(n4466), .IN5(
        n4814), .Q(n4805) );
  AO21X1 U4013 ( .IN1(N3708), .IN2(n4468), .IN3(n4469), .Q(n4814) );
  AO221X1 U4014 ( .IN1(N3811), .IN2(n4474), .IN3(N3744), .IN4(n4473), .IN5(
        n4815), .Q(n4804) );
  AO22X1 U4015 ( .IN1(N1201), .IN2(n4505), .IN3(N1233), .IN4(n4471), .Q(n4815)
         );
  MUX21X1 U4016 ( .IN1(n3831), .IN2(n4816), .S(n4438), .Q(n3471) );
  MUX21X1 U4017 ( .IN1(data_address[21]), .IN2(n4816), .S(n4439), .Q(n3470) );
  AO222X1 U4018 ( .IN1(n4434), .IN2(n293), .IN3(N1234), .IN4(n4435), .IN5(
        n4436), .IN6(SP[21]), .Q(n3469) );
  AO222X1 U4019 ( .IN1(n4440), .IN2(n3831), .IN3(n4441), .IN4(n4816), .IN5(
        n4442), .IN6(n3895), .Q(n3468) );
  OR4X1 U4020 ( .IN1(n4817), .IN2(n4818), .IN3(n4819), .IN4(n4820), .Q(n4816)
         );
  AO221X1 U4021 ( .IN1(n4454), .IN2(n4808), .IN3(n4463), .IN4(n4821), .IN5(
        n4822), .Q(n4820) );
  AO22X1 U4022 ( .IN1(N1169), .IN2(n4470), .IN3(n293), .IN4(n4457), .Q(n4822)
         );
  AO221X1 U4023 ( .IN1(n4452), .IN2(n4785), .IN3(n4459), .IN4(n4823), .IN5(
        n4824), .Q(n4819) );
  AO222X1 U4024 ( .IN1(n4449), .IN2(n4795), .IN3(n4825), .IN4(n4462), .IN5(
        n4447), .IN6(n4771), .Q(n4824) );
  AO222X1 U4025 ( .IN1(n4826), .IN2(n4827), .IN3(n4808), .IN4(n4761), .IN5(
        n4828), .IN6(n4829), .Q(n4771) );
  NOR2X0 U4026 ( .IN1(n3073), .IN2(n3020), .QN(n4825) );
  AO221X1 U4027 ( .IN1(n4758), .IN2(n4812), .IN3(n4830), .IN4(n4761), .IN5(
        n4794), .Q(n4795) );
  AO222X1 U4028 ( .IN1(n4797), .IN2(n4813), .IN3(n4753), .IN4(n4799), .IN5(
        n4831), .IN6(n4720), .Q(n4794) );
  AO222X1 U4029 ( .IN1(n4832), .IN2(n4833), .IN3(n4834), .IN4(n4835), .IN5(
        n4836), .IN6(n4837), .Q(n4799) );
  AO221X1 U4030 ( .IN1(N3577), .IN2(n4465), .IN3(N3848), .IN4(n4466), .IN5(
        n4838), .Q(n4818) );
  AO21X1 U4031 ( .IN1(N3709), .IN2(n4468), .IN3(n4469), .Q(n4838) );
  AO221X1 U4032 ( .IN1(N3812), .IN2(n4474), .IN3(N3745), .IN4(n4473), .IN5(
        n4839), .Q(n4817) );
  AO22X1 U4033 ( .IN1(N1202), .IN2(n4505), .IN3(N1234), .IN4(n4471), .Q(n4839)
         );
  MUX21X1 U4034 ( .IN1(n3832), .IN2(n4840), .S(n4438), .Q(n3467) );
  MUX21X1 U4035 ( .IN1(data_address[22]), .IN2(n4840), .S(n4439), .Q(n3466) );
  AO222X1 U4036 ( .IN1(n4434), .IN2(n292), .IN3(N1235), .IN4(n4435), .IN5(
        n4436), .IN6(SP[22]), .Q(n3465) );
  AO222X1 U4037 ( .IN1(n4440), .IN2(n3832), .IN3(n4441), .IN4(n4840), .IN5(
        n4442), .IN6(n3894), .Q(n3464) );
  OR4X1 U4038 ( .IN1(n4841), .IN2(n4842), .IN3(n4843), .IN4(n4844), .Q(n4840)
         );
  AO221X1 U4039 ( .IN1(n4454), .IN2(n4821), .IN3(n4463), .IN4(n4845), .IN5(
        n4846), .Q(n4844) );
  AO22X1 U4040 ( .IN1(N1170), .IN2(n4470), .IN3(n292), .IN4(n4457), .Q(n4846)
         );
  AO221X1 U4041 ( .IN1(n4452), .IN2(n4808), .IN3(n4459), .IN4(n4847), .IN5(
        n4848), .Q(n4843) );
  AO222X1 U4042 ( .IN1(n4447), .IN2(n4785), .IN3(n4849), .IN4(n4462), .IN5(
        n4449), .IN6(n4823), .Q(n4848) );
  AO221X1 U4043 ( .IN1(n4850), .IN2(n4761), .IN3(n4851), .IN4(n4691), .IN5(
        n4852), .Q(n4823) );
  AO22X1 U4044 ( .IN1(n4758), .IN2(n4830), .IN3(n4762), .IN4(n4812), .Q(n4852)
         );
  AO222X1 U4045 ( .IN1(n4797), .IN2(n4831), .IN3(n4753), .IN4(n4813), .IN5(
        n4853), .IN6(n4720), .Q(n4812) );
  AO222X1 U4046 ( .IN1(n4834), .IN2(n4854), .IN3(n4832), .IN4(n4835), .IN5(
        n4836), .IN6(n4833), .Q(n4813) );
  NOR2X0 U4047 ( .IN1(n3072), .IN2(n3018), .QN(n4849) );
  AO222X1 U4048 ( .IN1(n4821), .IN2(n4761), .IN3(n4828), .IN4(n4808), .IN5(
        n4826), .IN6(n4829), .Q(n4785) );
  AO221X1 U4049 ( .IN1(N3578), .IN2(n4465), .IN3(N3849), .IN4(n4466), .IN5(
        n4855), .Q(n4842) );
  AO21X1 U4050 ( .IN1(N3710), .IN2(n4468), .IN3(n4469), .Q(n4855) );
  AO221X1 U4051 ( .IN1(N3813), .IN2(n4474), .IN3(N3746), .IN4(n4473), .IN5(
        n4856), .Q(n4841) );
  AO22X1 U4052 ( .IN1(N1203), .IN2(n4505), .IN3(N1235), .IN4(n4471), .Q(n4856)
         );
  MUX21X1 U4053 ( .IN1(n3833), .IN2(n4857), .S(n4438), .Q(n3463) );
  MUX21X1 U4054 ( .IN1(data_address[23]), .IN2(n4857), .S(n4439), .Q(n3462) );
  AO222X1 U4055 ( .IN1(n4434), .IN2(n291), .IN3(N1236), .IN4(n4435), .IN5(
        n4436), .IN6(SP[23]), .Q(n3461) );
  AO222X1 U4056 ( .IN1(n4440), .IN2(n3833), .IN3(n4441), .IN4(n4857), .IN5(
        n4442), .IN6(n3893), .Q(n3460) );
  OR4X1 U4057 ( .IN1(n4858), .IN2(n4859), .IN3(n4860), .IN4(n4861), .Q(n4857)
         );
  AO221X1 U4058 ( .IN1(n4454), .IN2(n4845), .IN3(n4459), .IN4(n4862), .IN5(
        n4863), .Q(n4861) );
  AO22X1 U4059 ( .IN1(N1171), .IN2(n4470), .IN3(n291), .IN4(n4457), .Q(n4863)
         );
  AO221X1 U4060 ( .IN1(n4449), .IN2(n4847), .IN3(n4452), .IN4(n4821), .IN5(
        n4864), .Q(n4860) );
  AO22X1 U4061 ( .IN1(n4447), .IN2(n4808), .IN3(n4865), .IN4(n4462), .Q(n4864)
         );
  NOR2X0 U4062 ( .IN1(n3071), .IN2(n3016), .QN(n4865) );
  AO222X1 U4063 ( .IN1(n4866), .IN2(n4867), .IN3(n4868), .IN4(n4845), .IN5(
        n4869), .IN6(n4870), .Q(n4808) );
  AO221X1 U4064 ( .IN1(n4871), .IN2(n4761), .IN3(n4872), .IN4(n4691), .IN5(
        n4873), .Q(n4847) );
  AO22X1 U4065 ( .IN1(n4758), .IN2(n4850), .IN3(n4762), .IN4(n4830), .Q(n4873)
         );
  AO222X1 U4066 ( .IN1(n4797), .IN2(n4853), .IN3(n4753), .IN4(n4831), .IN5(
        n4874), .IN6(n4720), .Q(n4830) );
  AO221X1 U4067 ( .IN1(n4832), .IN2(n4854), .IN3(n4834), .IN4(n4875), .IN5(
        n4835), .Q(n4831) );
  AO222X1 U4068 ( .IN1(n4876), .IN2(n4877), .IN3(n4878), .IN4(n4879), .IN5(
        n4880), .IN6(n4881), .Q(n4835) );
  AO221X1 U4069 ( .IN1(N3579), .IN2(n4465), .IN3(N3850), .IN4(n4466), .IN5(
        n4882), .Q(n4859) );
  AO21X1 U4070 ( .IN1(N3711), .IN2(n4468), .IN3(n4883), .Q(n4882) );
  AO221X1 U4071 ( .IN1(N3814), .IN2(n4474), .IN3(N3747), .IN4(n4473), .IN5(
        n4884), .Q(n4858) );
  AO22X1 U4072 ( .IN1(N1204), .IN2(n4505), .IN3(N1236), .IN4(n4471), .Q(n4884)
         );
  MUX21X1 U4073 ( .IN1(n3834), .IN2(n4885), .S(n4438), .Q(n3459) );
  MUX21X1 U4074 ( .IN1(data_address[24]), .IN2(n4885), .S(n4439), .Q(n3458) );
  AO222X1 U4075 ( .IN1(n4434), .IN2(n290), .IN3(N1237), .IN4(n4435), .IN5(
        n4436), .IN6(SP[24]), .Q(n3457) );
  AO222X1 U4076 ( .IN1(n4440), .IN2(n3834), .IN3(n4441), .IN4(n4885), .IN5(
        n4442), .IN6(n3892), .Q(n3456) );
  OR4X1 U4077 ( .IN1(n4886), .IN2(n4887), .IN3(n4888), .IN4(n4889), .Q(n4885)
         );
  AO221X1 U4078 ( .IN1(n4459), .IN2(n4890), .IN3(n290), .IN4(n4457), .IN5(
        n4891), .Q(n4889) );
  AO222X1 U4079 ( .IN1(n4454), .IN2(n4892), .IN3(n4452), .IN4(n4845), .IN5(
        n4893), .IN6(n4862), .Q(n4891) );
  AO221X1 U4080 ( .IN1(n4447), .IN2(n4821), .IN3(n4894), .IN4(n4872), .IN5(
        n4895), .Q(n4888) );
  AO222X1 U4081 ( .IN1(n4463), .IN2(n4896), .IN3(n4897), .IN4(n4462), .IN5(
        n4898), .IN6(n4899), .Q(n4895) );
  AO222X1 U4082 ( .IN1(n4621), .IN2(n4872), .IN3(n4624), .IN4(n4851), .IN5(
        n4862), .IN6(n4591), .Q(n4899) );
  AO221X1 U4083 ( .IN1(n4900), .IN2(n4761), .IN3(n4724), .IN4(n4872), .IN5(
        n4901), .Q(n4851) );
  AO22X1 U4084 ( .IN1(n4758), .IN2(n4871), .IN3(n4762), .IN4(n4850), .Q(n4901)
         );
  AO222X1 U4085 ( .IN1(n4797), .IN2(n4874), .IN3(n4753), .IN4(n4853), .IN5(
        n4902), .IN6(n4720), .Q(n4850) );
  AO21X1 U4086 ( .IN1(n4832), .IN2(n4875), .IN3(n4854), .Q(n4853) );
  AO222X1 U4087 ( .IN1(n4903), .IN2(n4879), .IN3(n4876), .IN4(n4878), .IN5(
        n4880), .IN6(n4877), .Q(n4854) );
  NOR2X0 U4088 ( .IN1(n3070), .IN2(n3014), .QN(n4897) );
  AO222X1 U4089 ( .IN1(n4868), .IN2(n4904), .IN3(n4869), .IN4(n4845), .IN5(
        n4866), .IN6(n4870), .Q(n4821) );
  AO221X1 U4090 ( .IN1(N3580), .IN2(n4465), .IN3(N3851), .IN4(n4466), .IN5(
        n4905), .Q(n4887) );
  AO21X1 U4091 ( .IN1(N3712), .IN2(n4468), .IN3(n4469), .Q(n4905) );
  AO221X1 U4092 ( .IN1(N3815), .IN2(n4474), .IN3(N3748), .IN4(n4473), .IN5(
        n4906), .Q(n4886) );
  AO222X1 U4093 ( .IN1(N1237), .IN2(n4471), .IN3(N1172), .IN4(n4470), .IN5(
        N1205), .IN6(n4505), .Q(n4906) );
  MUX21X1 U4094 ( .IN1(n3835), .IN2(n4907), .S(n4438), .Q(n3455) );
  MUX21X1 U4095 ( .IN1(data_address[25]), .IN2(n4907), .S(n4439), .Q(n3454) );
  AO222X1 U4096 ( .IN1(n4434), .IN2(n289), .IN3(N1238), .IN4(n4435), .IN5(
        n4436), .IN6(SP[25]), .Q(n3453) );
  AO222X1 U4097 ( .IN1(n4440), .IN2(n3835), .IN3(n4441), .IN4(n4907), .IN5(
        n4442), .IN6(n3891), .Q(n3452) );
  OR4X1 U4098 ( .IN1(n4908), .IN2(n4909), .IN3(n4910), .IN4(n4911), .Q(n4907)
         );
  AO221X1 U4099 ( .IN1(n4893), .IN2(n4890), .IN3(n4454), .IN4(n4896), .IN5(
        n4912), .Q(n4911) );
  AO22X1 U4100 ( .IN1(n289), .IN2(n4457), .IN3(n4459), .IN4(n4913), .Q(n4912)
         );
  AO221X1 U4101 ( .IN1(n4452), .IN2(n4892), .IN3(n4894), .IN4(n4862), .IN5(
        n4914), .Q(n4910) );
  AO222X1 U4102 ( .IN1(n4898), .IN2(n4872), .IN3(n4915), .IN4(n4462), .IN5(
        n4447), .IN6(n4845), .Q(n4914) );
  AO222X1 U4103 ( .IN1(n4916), .IN2(n4917), .IN3(n4918), .IN4(n4919), .IN5(
        n4920), .IN6(n4921), .Q(n4845) );
  NOR2X0 U4104 ( .IN1(n3069), .IN2(n3012), .QN(n4915) );
  AO221X1 U4105 ( .IN1(n4758), .IN2(n4900), .IN3(n4922), .IN4(n4761), .IN5(
        n4871), .Q(n4872) );
  AO222X1 U4106 ( .IN1(n4797), .IN2(n4902), .IN3(n4753), .IN4(n4874), .IN5(
        n4923), .IN6(n4720), .Q(n4871) );
  AO21X1 U4107 ( .IN1(n4832), .IN2(n4924), .IN3(n4875), .Q(n4874) );
  AO221X1 U4108 ( .IN1(n4876), .IN2(n4903), .IN3(n4925), .IN4(n4879), .IN5(
        n4878), .Q(n4875) );
  AO222X1 U4109 ( .IN1(n4926), .IN2(n4927), .IN3(n4928), .IN4(n4929), .IN5(
        n4930), .IN6(n4931), .Q(n4878) );
  AO221X1 U4110 ( .IN1(N3581), .IN2(n4465), .IN3(N3852), .IN4(n4466), .IN5(
        n4932), .Q(n4909) );
  AO21X1 U4111 ( .IN1(N3713), .IN2(n4468), .IN3(n4883), .Q(n4932) );
  AO21X1 U4112 ( .IN1(n4463), .IN2(n4892), .IN3(n4469), .Q(n4883) );
  AO221X1 U4113 ( .IN1(N3816), .IN2(n4474), .IN3(N3749), .IN4(n4473), .IN5(
        n4933), .Q(n4908) );
  AO222X1 U4114 ( .IN1(N1238), .IN2(n4471), .IN3(N1173), .IN4(n4470), .IN5(
        N1206), .IN6(n4505), .Q(n4933) );
  MUX21X1 U4115 ( .IN1(n3836), .IN2(n4934), .S(n4438), .Q(n3451) );
  MUX21X1 U4116 ( .IN1(data_address[26]), .IN2(n4934), .S(n4439), .Q(n3450) );
  AO222X1 U4117 ( .IN1(n4434), .IN2(n288), .IN3(N1239), .IN4(n4435), .IN5(
        n4436), .IN6(SP[26]), .Q(n3449) );
  AO222X1 U4118 ( .IN1(n4440), .IN2(n3836), .IN3(n4441), .IN4(n4934), .IN5(
        n4442), .IN6(n3890), .Q(n3448) );
  OR4X1 U4119 ( .IN1(n4935), .IN2(n4936), .IN3(n4937), .IN4(n4938), .Q(n4934)
         );
  AO221X1 U4120 ( .IN1(n4893), .IN2(n4913), .IN3(n4459), .IN4(n4939), .IN5(
        n4940), .Q(n4938) );
  AO22X1 U4121 ( .IN1(N1174), .IN2(n4470), .IN3(n288), .IN4(n4457), .Q(n4940)
         );
  AO221X1 U4122 ( .IN1(n4894), .IN2(n4890), .IN3(n4463), .IN4(n4896), .IN5(
        n4941), .Q(n4937) );
  AO222X1 U4123 ( .IN1(n4942), .IN2(n4892), .IN3(n4943), .IN4(n4462), .IN5(
        n4898), .IN6(n4862), .Q(n4941) );
  AO222X1 U4124 ( .IN1(n4758), .IN2(n4922), .IN3(n4762), .IN4(n4900), .IN5(
        n4913), .IN6(n4761), .Q(n4862) );
  AO222X1 U4125 ( .IN1(n4797), .IN2(n4923), .IN3(n4753), .IN4(n4902), .IN5(
        n4944), .IN6(n4720), .Q(n4900) );
  AO21X1 U4126 ( .IN1(n4832), .IN2(n4925), .IN3(n4924), .Q(n4902) );
  AO21X1 U4127 ( .IN1(n4876), .IN2(n4925), .IN3(n4903), .Q(n4924) );
  AO222X1 U4128 ( .IN1(n4928), .IN2(n4945), .IN3(n4926), .IN4(n4929), .IN5(
        n4930), .IN6(n4927), .Q(n4903) );
  NOR2X0 U4129 ( .IN1(n3068), .IN2(n3010), .QN(n4943) );
  AO222X1 U4130 ( .IN1(n4792), .IN2(n4946), .IN3(n4789), .IN4(n4947), .IN5(
        n4948), .IN6(n4791), .Q(n4892) );
  AO221X1 U4131 ( .IN1(n4828), .IN2(n4949), .IN3(n4948), .IN4(n4761), .IN5(
        n4904), .Q(n4947) );
  AO222X1 U4132 ( .IN1(n4950), .IN2(n4919), .IN3(n4920), .IN4(n4918), .IN5(
        n4916), .IN6(n4921), .Q(n4904) );
  AO221X1 U4133 ( .IN1(N3582), .IN2(n4465), .IN3(N3853), .IN4(n4466), .IN5(
        n4951), .Q(n4936) );
  AO21X1 U4134 ( .IN1(N3714), .IN2(n4468), .IN3(n4469), .Q(n4951) );
  AO221X1 U4135 ( .IN1(N3817), .IN2(n4474), .IN3(N3750), .IN4(n4473), .IN5(
        n4952), .Q(n4935) );
  AO22X1 U4136 ( .IN1(N1207), .IN2(n4505), .IN3(N1239), .IN4(n4471), .Q(n4952)
         );
  MUX21X1 U4137 ( .IN1(n3837), .IN2(n4953), .S(n4438), .Q(n3447) );
  MUX21X1 U4138 ( .IN1(data_address[27]), .IN2(n4953), .S(n4439), .Q(n3446) );
  AO222X1 U4139 ( .IN1(n4434), .IN2(n287), .IN3(N1240), .IN4(n4435), .IN5(
        n4436), .IN6(SP[27]), .Q(n3445) );
  AO222X1 U4140 ( .IN1(n4440), .IN2(n3837), .IN3(n4441), .IN4(n4953), .IN5(
        n4442), .IN6(n3889), .Q(n3444) );
  OR4X1 U4141 ( .IN1(n4954), .IN2(n4955), .IN3(n4956), .IN4(n4957), .Q(n4953)
         );
  AO221X1 U4142 ( .IN1(n4894), .IN2(n4913), .IN3(n4893), .IN4(n4939), .IN5(
        n4958), .Q(n4957) );
  AO22X1 U4143 ( .IN1(N1175), .IN2(n4470), .IN3(n287), .IN4(n4457), .Q(n4958)
         );
  AO221X1 U4144 ( .IN1(n4898), .IN2(n4890), .IN3(n4942), .IN4(n4896), .IN5(
        n4959), .Q(n4956) );
  AO22X1 U4145 ( .IN1(n4463), .IN2(n4948), .IN3(n4960), .IN4(n4462), .Q(n4959)
         );
  NOR2X0 U4146 ( .IN1(n3067), .IN2(n3008), .QN(n4960) );
  AO222X1 U4147 ( .IN1(n4792), .IN2(n4948), .IN3(n4789), .IN4(n4946), .IN5(
        n4961), .IN6(n4791), .Q(n4896) );
  AO21X1 U4148 ( .IN1(n4828), .IN2(n4948), .IN3(n4949), .Q(n4946) );
  AO221X1 U4149 ( .IN1(n4920), .IN2(n4950), .IN3(n4962), .IN4(n4919), .IN5(
        n4918), .Q(n4949) );
  AO222X1 U4150 ( .IN1(n4727), .IN2(n4963), .IN3(n4964), .IN4(n4965), .IN5(
        n4966), .IN6(n4967), .Q(n4918) );
  AO222X1 U4151 ( .IN1(n4758), .IN2(n4913), .IN3(n4762), .IN4(n4922), .IN5(
        n4939), .IN6(n4761), .Q(n4890) );
  AO222X1 U4152 ( .IN1(n4797), .IN2(n4944), .IN3(n4753), .IN4(n4923), .IN5(
        n4968), .IN6(n4720), .Q(n4922) );
  AO21X1 U4153 ( .IN1(n4832), .IN2(n4944), .IN3(n4925), .Q(n4923) );
  AO222X1 U4154 ( .IN1(n4926), .IN2(n4945), .IN3(n4930), .IN4(n4929), .IN5(
        n4928), .IN6(n4969), .Q(n4925) );
  AO222X1 U4155 ( .IN1(n4970), .IN2(n4971), .IN3(n4972), .IN4(n4973), .IN5(
        n4974), .IN6(n4975), .Q(n4929) );
  AO221X1 U4156 ( .IN1(N3583), .IN2(n4465), .IN3(N3854), .IN4(n4466), .IN5(
        n4976), .Q(n4955) );
  AO21X1 U4157 ( .IN1(N3715), .IN2(n4468), .IN3(n4977), .Q(n4976) );
  AO221X1 U4158 ( .IN1(N3818), .IN2(n4474), .IN3(N3751), .IN4(n4473), .IN5(
        n4978), .Q(n4954) );
  AO22X1 U4159 ( .IN1(N1208), .IN2(n4505), .IN3(N1240), .IN4(n4471), .Q(n4978)
         );
  MUX21X1 U4160 ( .IN1(n3838), .IN2(n4979), .S(n4438), .Q(n3443) );
  MUX21X1 U4161 ( .IN1(data_address[28]), .IN2(n4979), .S(n4439), .Q(n3442) );
  AO222X1 U4162 ( .IN1(n4434), .IN2(n286), .IN3(N1241), .IN4(n4435), .IN5(
        n4436), .IN6(SP[28]), .Q(n3441) );
  AO222X1 U4163 ( .IN1(n4440), .IN2(n3838), .IN3(n4441), .IN4(n4979), .IN5(
        n4442), .IN6(n3888), .Q(n3440) );
  OR4X1 U4164 ( .IN1(n4980), .IN2(n4981), .IN3(n4982), .IN4(n4983), .Q(n4979)
         );
  AO221X1 U4165 ( .IN1(n4894), .IN2(n4939), .IN3(n286), .IN4(n4457), .IN5(
        n4984), .Q(n4983) );
  AO22X1 U4166 ( .IN1(N1241), .IN2(n4471), .IN3(N1176), .IN4(n4470), .Q(n4984)
         );
  AO221X1 U4167 ( .IN1(n4898), .IN2(n4913), .IN3(n4463), .IN4(n4961), .IN5(
        n4985), .Q(n4982) );
  AO22X1 U4168 ( .IN1(n4942), .IN2(n4948), .IN3(n4986), .IN4(n4462), .Q(n4985)
         );
  NOR2X0 U4169 ( .IN1(n3066), .IN2(n3006), .QN(n4986) );
  AO221X1 U4170 ( .IN1(n4920), .IN2(n4962), .IN3(n4987), .IN4(n4919), .IN5(
        n4950), .Q(n4948) );
  AO222X1 U4171 ( .IN1(n4987), .IN2(n4965), .IN3(n4966), .IN4(n4964), .IN5(
        n4727), .IN6(n4967), .Q(n4950) );
  AO222X1 U4172 ( .IN1(n4797), .IN2(n4968), .IN3(n4753), .IN4(n4944), .IN5(
        n4988), .IN6(n4720), .Q(n4913) );
  AO222X1 U4173 ( .IN1(n4926), .IN2(n4969), .IN3(n4930), .IN4(n4945), .IN5(
        n4928), .IN6(n4988), .Q(n4944) );
  AO222X1 U4174 ( .IN1(n4988), .IN2(n4973), .IN3(n4970), .IN4(n4972), .IN5(
        n4974), .IN6(n4971), .Q(n4945) );
  AO221X1 U4175 ( .IN1(N3855), .IN2(n4466), .IN3(N3716), .IN4(n4468), .IN5(
        n4989), .Q(n4981) );
  AO221X1 U4176 ( .IN1(N3752), .IN2(n4473), .IN3(N3584), .IN4(n4465), .IN5(
        n4990), .Q(n4980) );
  AO22X1 U4177 ( .IN1(N3819), .IN2(n4474), .IN3(N1209), .IN4(n4505), .Q(n4990)
         );
  MUX21X1 U4178 ( .IN1(n3839), .IN2(n4991), .S(n4438), .Q(n3439) );
  MUX21X1 U4179 ( .IN1(data_address[29]), .IN2(n4991), .S(n4439), .Q(n3438) );
  AO222X1 U4180 ( .IN1(n4434), .IN2(n285), .IN3(N1242), .IN4(n4435), .IN5(
        n4436), .IN6(SP[29]), .Q(n3437) );
  AO222X1 U4181 ( .IN1(n4440), .IN2(n3839), .IN3(n4441), .IN4(n4991), .IN5(
        n4442), .IN6(n3887), .Q(n3436) );
  OR4X1 U4182 ( .IN1(n4992), .IN2(n4993), .IN3(n4994), .IN4(n4995), .Q(n4991)
         );
  AO221X1 U4183 ( .IN1(N1177), .IN2(n4470), .IN3(N1242), .IN4(n4471), .IN5(
        n4996), .Q(n4995) );
  AO22X1 U4184 ( .IN1(n4463), .IN2(n4357), .IN3(n285), .IN4(n4457), .Q(n4996)
         );
  AO221X1 U4185 ( .IN1(n4997), .IN2(n4462), .IN3(n4942), .IN4(n4961), .IN5(
        n4998), .Q(n4994) );
  AO22X1 U4186 ( .IN1(n4894), .IN2(n4296), .IN3(n4898), .IN4(n4939), .Q(n4998)
         );
  AO222X1 U4187 ( .IN1(n4797), .IN2(n4988), .IN3(n4753), .IN4(n4968), .IN5(
        n4720), .IN6(n4296), .Q(n4939) );
  AO222X1 U4188 ( .IN1(n4988), .IN2(n4926), .IN3(n4930), .IN4(n4969), .IN5(
        n4928), .IN6(n4296), .Q(n4968) );
  AO221X1 U4189 ( .IN1(n4970), .IN2(n4988), .IN3(n4973), .IN4(n4296), .IN5(
        n4972), .Q(n4969) );
  AO22X1 U4190 ( .IN1(n4999), .IN2(n4295), .IN3(n5000), .IN4(n4296), .Q(n4972)
         );
  NOR2X0 U4191 ( .IN1(n5001), .IN2(n5725), .QN(n4988) );
  AO222X1 U4192 ( .IN1(n4987), .IN2(n4869), .IN3(n4866), .IN4(n4962), .IN5(
        n4868), .IN6(n4357), .Q(n4961) );
  AO21X1 U4193 ( .IN1(n4966), .IN2(n4987), .IN3(n4964), .Q(n4962) );
  AO222X1 U4194 ( .IN1(n5002), .IN2(n4357), .IN3(n5003), .IN4(n4355), .IN5(
        n5004), .IN6(n4356), .Q(n4964) );
  NOR2X0 U4195 ( .IN1(n3065), .IN2(n3004), .QN(n4997) );
  AO221X1 U4196 ( .IN1(N3856), .IN2(n4466), .IN3(N3717), .IN4(n4468), .IN5(
        n4989), .Q(n4993) );
  AO21X1 U4197 ( .IN1(n4893), .IN2(n4296), .IN3(n4977), .Q(n4989) );
  AO21X1 U4198 ( .IN1(n4459), .IN2(n4296), .IN3(n4469), .Q(n4977) );
  AO221X1 U4199 ( .IN1(N3753), .IN2(n4473), .IN3(N3585), .IN4(n4465), .IN5(
        n5005), .Q(n4992) );
  AO22X1 U4200 ( .IN1(N3820), .IN2(n4474), .IN3(N1210), .IN4(n4505), .Q(n5005)
         );
  MUX21X1 U4201 ( .IN1(n3840), .IN2(n5006), .S(n4438), .Q(n3435) );
  MUX21X1 U4202 ( .IN1(data_address[30]), .IN2(n5006), .S(n4439), .Q(n3434) );
  AO222X1 U4203 ( .IN1(n4434), .IN2(n284), .IN3(N1243), .IN4(n4435), .IN5(
        n4436), .IN6(SP[30]), .Q(n3433) );
  NOR2X0 U4204 ( .IN1(n4436), .IN2(n5724), .QN(n4435) );
  NOR2X0 U4205 ( .IN1(n4436), .IN2(n3843), .QN(n4434) );
  NAND2X0 U4206 ( .IN1(n5007), .IN2(n4254), .QN(n4436) );
  MUX21X1 U4207 ( .IN1(n5008), .IN2(n4505), .S(n5722), .Q(n5007) );
  AO222X1 U4208 ( .IN1(n4440), .IN2(n3840), .IN3(n4441), .IN4(n5006), .IN5(
        n4442), .IN6(n3886), .Q(n3432) );
  OR4X1 U4209 ( .IN1(n5009), .IN2(n5010), .IN3(n5011), .IN4(n5012), .Q(n5006)
         );
  AO222X1 U4210 ( .IN1(N1178), .IN2(n4470), .IN3(n284), .IN4(n4457), .IN5(
        N1243), .IN6(n4471), .Q(n5012) );
  NAND3X0 U4211 ( .IN1(n5013), .IN2(n5014), .IN3(n5015), .QN(n5011) );
  AOI22X1 U4212 ( .IN1(n4357), .IN2(n5016), .IN3(n4987), .IN4(n4447), .QN(
        n5015) );
  MUX21X1 U4213 ( .IN1(n4357), .IN2(n4356), .S(n5003), .Q(n4987) );
  AO21X1 U4214 ( .IN1(n5017), .IN2(n4942), .IN3(n4463), .Q(n5016) );
  NAND3X0 U4215 ( .IN1(n4356), .IN2(n4295), .IN3(n4462), .QN(n5013) );
  AO221X1 U4216 ( .IN1(N3857), .IN2(n4466), .IN3(N3718), .IN4(n4468), .IN5(
        n4469), .Q(n5010) );
  AO221X1 U4217 ( .IN1(N3754), .IN2(n4473), .IN3(N3586), .IN4(n4465), .IN5(
        n5018), .Q(n5009) );
  AO22X1 U4218 ( .IN1(N3821), .IN2(n4474), .IN3(N1211), .IN4(n4505), .Q(n5018)
         );
  MUX21X1 U4219 ( .IN1(n3841), .IN2(n4416), .S(n4438), .Q(n3431) );
  MUX21X1 U4220 ( .IN1(data_address[31]), .IN2(n4416), .S(n4439), .Q(n3430) );
  AO222X1 U4221 ( .IN1(n4440), .IN2(n3841), .IN3(n4441), .IN4(n4416), .IN5(
        n4442), .IN6(n3885), .Q(n3429) );
  OR4X1 U4222 ( .IN1(n5021), .IN2(n5022), .IN3(n5023), .IN4(n5024), .Q(n4416)
         );
  AO222X1 U4223 ( .IN1(N1212), .IN2(n4505), .IN3(N1244), .IN4(n4471), .IN5(
        N3719), .IN6(n4468), .Q(n5024) );
  AO221X1 U4224 ( .IN1(N3822), .IN2(n4474), .IN3(N3587), .IN4(n4465), .IN5(
        n5025), .Q(n5023) );
  NAND2X0 U4225 ( .IN1(n5026), .IN2(n5014), .QN(n5025) );
  NAND3X0 U4226 ( .IN1(n4357), .IN2(n4296), .IN3(n4462), .QN(n5026) );
  NOR3X0 U4227 ( .IN1(n3804), .IN2(n5723), .IN3(n3807), .QN(n4462) );
  AO222X1 U4228 ( .IN1(n5027), .IN2(n4357), .IN3(n283), .IN4(n4457), .IN5(
        N3755), .IN6(n4473), .Q(n5022) );
  AO221X1 U4229 ( .IN1(n5028), .IN2(n5029), .IN3(n5030), .IN4(n5721), .IN5(
        n5031), .Q(n4457) );
  NOR2X0 U4230 ( .IN1(n5724), .IN2(n5032), .QN(n5028) );
  AO221X1 U4231 ( .IN1(N1179), .IN2(n4470), .IN3(N3858), .IN4(n4466), .IN5(
        n5033), .Q(n5021) );
  AND2X1 U4232 ( .IN1(n5034), .IN2(n5035), .Q(n4441) );
  AND2X1 U4233 ( .IN1(n5019), .IN2(n5034), .Q(n4440) );
  NOR2X0 U4234 ( .IN1(n4442), .IN2(n5036), .QN(n5034) );
  AND4X1 U4235 ( .IN1(n4418), .IN2(n4423), .IN3(n5037), .IN4(n5038), .Q(n5036)
         );
  OA221X1 U4236 ( .IN1(n4429), .IN2(n5039), .IN3(n5040), .IN4(n3807), .IN5(
        n5041), .Q(n5038) );
  OA22X1 U4237 ( .IN1(n5042), .IN2(n5043), .IN3(n4417), .IN4(n5044), .Q(n5041)
         );
  OA21X1 U4238 ( .IN1(n3804), .IN2(n4582), .IN3(n5045), .Q(n5040) );
  MUX21X1 U4239 ( .IN1(n5046), .IN2(n5047), .S(\r150/A[3] ), .Q(n5037) );
  NAND2X0 U4240 ( .IN1(n4427), .IN2(n3843), .QN(n5047) );
  NAND2X0 U4241 ( .IN1(n5721), .IN2(n5048), .QN(n5046) );
  OA22X1 U4242 ( .IN1(n5049), .IN2(n4428), .IN3(n5722), .IN4(n5050), .Q(n4423)
         );
  AOI21X1 U4243 ( .IN1(n4406), .IN2(n4407), .IN3(n5008), .QN(n5050) );
  NOR2X0 U4244 ( .IN1(n3803), .IN2(n4433), .QN(n5008) );
  AND2X1 U4245 ( .IN1(n4404), .IN2(n5051), .Q(n4418) );
  NAND3X0 U4246 ( .IN1(n5721), .IN2(n5723), .IN3(n4410), .QN(n5051) );
  NAND3X0 U4247 ( .IN1(n4409), .IN2(n3803), .IN3(n5052), .QN(n4404) );
  NAND2X0 U4248 ( .IN1(n4254), .IN2(n5020), .QN(n4442) );
  NAND4X0 U4249 ( .IN1(n5053), .IN2(n5054), .IN3(n5045), .IN4(n5049), .QN(
        n5020) );
  NAND3X0 U4250 ( .IN1(n4429), .IN2(n3804), .IN3(n5048), .QN(n5049) );
  NAND2X0 U4251 ( .IN1(n4406), .IN2(n5723), .QN(n5054) );
  MUX21X1 U4252 ( .IN1(n3804), .IN2(n5048), .S(n4428), .Q(n5053) );
  INVX0 U4253 ( .INP(n4400), .ZN(n4254) );
  INVX0 U4254 ( .INP(n5035), .ZN(n5019) );
  NAND3X0 U4255 ( .IN1(n5055), .IN2(n5056), .IN3(n5057), .QN(n5035) );
  AO21X1 U4256 ( .IN1(n4406), .IN2(n3805), .IN3(n3804), .Q(n5057) );
  MUX21X1 U4257 ( .IN1(n3847), .IN2(n4430), .S(n5058), .Q(n3428) );
  NOR2X0 U4258 ( .IN1(n4431), .IN2(n4400), .QN(n5058) );
  NAND2X0 U4259 ( .IN1(reset_n), .IN2(n5711), .QN(n4400) );
  AND4X1 U4260 ( .IN1(n5055), .IN2(n5043), .IN3(n5059), .IN4(n5060), .Q(n4431)
         );
  NAND2X0 U4261 ( .IN1(n4420), .IN2(n5032), .QN(n5060) );
  NOR2X0 U4262 ( .IN1(n4425), .IN2(n5052), .QN(n5059) );
  AND2X1 U4263 ( .IN1(n5722), .IN2(n4407), .Q(n5052) );
  NAND2X0 U4264 ( .IN1(n3805), .IN2(n4429), .QN(n5043) );
  NAND2X0 U4265 ( .IN1(n3804), .IN2(n4433), .QN(n5055) );
  NAND2X0 U4266 ( .IN1(n4407), .IN2(n4428), .QN(n4433) );
  OR4X1 U4267 ( .IN1(n5061), .IN2(n5062), .IN3(n5063), .IN4(n5064), .Q(n4430)
         );
  AO221X1 U4268 ( .IN1(n4452), .IN2(n4448), .IN3(n4463), .IN4(n4455), .IN5(
        n5065), .Q(n5064) );
  AO22X1 U4269 ( .IN1(N1180), .IN2(n4470), .IN3(n4893), .IN4(n4490), .Q(n5065)
         );
  AND2X1 U4270 ( .IN1(n4449), .IN2(n4488), .Q(n4893) );
  OAI22X1 U4271 ( .IN1(n5722), .IN2(n5066), .IN3(n5056), .IN4(n5067), .QN(
        n4470) );
  MUX21X1 U4272 ( .IN1(n5068), .IN2(n3807), .S(n5723), .Q(n5067) );
  NAND2X0 U4273 ( .IN1(n5722), .IN2(n4428), .QN(n5068) );
  INVX0 U4274 ( .INP(n4409), .ZN(n4428) );
  NAND2X0 U4275 ( .IN1(n3844), .IN2(n3807), .QN(n4409) );
  OA21X1 U4276 ( .IN1(n5069), .IN2(n5032), .IN3(n5070), .Q(n5066) );
  NAND4X0 U4277 ( .IN1(n5721), .IN2(n5071), .IN3(n5072), .IN4(n5073), .QN(
        n5070) );
  NAND2X0 U4278 ( .IN1(n5029), .IN2(n5720), .QN(n5072) );
  INVX0 U4279 ( .INP(n5074), .ZN(n5029) );
  NAND2X0 U4280 ( .IN1(n5723), .IN2(n5075), .QN(n5071) );
  OA21X1 U4281 ( .IN1(n3843), .IN2(n5074), .IN3(n4582), .Q(n5069) );
  AO222X1 U4282 ( .IN1(n4518), .IN2(n4488), .IN3(n4517), .IN4(n4516), .IN5(
        n4515), .IN6(n5076), .Q(n4455) );
  AO222X1 U4283 ( .IN1(n4552), .IN2(n4522), .IN3(n4551), .IN4(n4550), .IN5(
        n4549), .IN6(n5077), .Q(n4518) );
  AO222X1 U4284 ( .IN1(n4593), .IN2(n4591), .IN3(n4592), .IN4(n4590), .IN5(
        n4589), .IN6(n5078), .Q(n4552) );
  AO222X1 U4285 ( .IN1(n4620), .IN2(n4618), .IN3(n4619), .IN4(n4617), .IN5(
        n4557), .IN6(n5079), .Q(n4593) );
  AO222X1 U4286 ( .IN1(n4653), .IN2(n4651), .IN3(n4652), .IN4(n4650), .IN5(
        n4649), .IN6(n5080), .Q(n4620) );
  AO222X1 U4287 ( .IN1(n4687), .IN2(n4685), .IN3(n4686), .IN4(n4684), .IN5(
        n4683), .IN6(n5081), .Q(n4653) );
  AO222X1 U4288 ( .IN1(n4722), .IN2(n4720), .IN3(n4721), .IN4(n4719), .IN5(
        n4718), .IN6(n5082), .Q(n4687) );
  AO222X1 U4289 ( .IN1(n4757), .IN2(n4755), .IN3(n4756), .IN4(n4754), .IN5(
        n4753), .IN6(n5083), .Q(n4722) );
  AO222X1 U4290 ( .IN1(n4793), .IN2(n4791), .IN3(n4792), .IN4(n4790), .IN5(
        n4789), .IN6(n5084), .Q(n4757) );
  AO222X1 U4291 ( .IN1(n4829), .IN2(n4761), .IN3(n4828), .IN4(n4827), .IN5(
        n4826), .IN6(n5085), .Q(n4793) );
  AO222X1 U4292 ( .IN1(n4868), .IN2(n4870), .IN3(n4869), .IN4(n4867), .IN5(
        n4866), .IN6(n5086), .Q(n4829) );
  AO222X1 U4293 ( .IN1(n4921), .IN2(n4919), .IN3(n4920), .IN4(n4917), .IN5(
        n4916), .IN6(n5087), .Q(n4870) );
  AO222X1 U4294 ( .IN1(n4967), .IN2(n4965), .IN3(n4966), .IN4(n4963), .IN5(
        n4727), .IN6(n5088), .Q(n4921) );
  AO222X1 U4295 ( .IN1(n5002), .IN2(n4356), .IN3(n5003), .IN4(n4354), .IN5(
        n5004), .IN6(n4355), .Q(n4967) );
  AND2X1 U4296 ( .IN1(n5089), .IN2(n5027), .Q(n4463) );
  AO222X1 U4297 ( .IN1(n4517), .IN2(n5090), .IN3(n5076), .IN4(n4488), .IN5(
        n4515), .IN6(n5091), .Q(n4448) );
  NOR3X0 U4298 ( .IN1(n4726), .IN2(n4523), .IN3(n5092), .QN(n4452) );
  AO221X1 U4299 ( .IN1(n4894), .IN2(n5093), .IN3(n4454), .IN4(n4453), .IN5(
        n5094), .Q(n5063) );
  AO222X1 U4300 ( .IN1(n4447), .IN2(n5095), .IN3(n4898), .IN4(n5096), .IN5(
        n282), .IN6(n5097), .Q(n5094) );
  AO221X1 U4301 ( .IN1(n5030), .IN2(n5722), .IN3(n4427), .IN4(n5048), .IN5(
        n5031), .Q(n5097) );
  AO221X1 U4302 ( .IN1(n4425), .IN2(n4427), .IN3(n4406), .IN4(n4407), .IN5(
        n5098), .Q(n5031) );
  INVX0 U4303 ( .INP(n5045), .ZN(n5098) );
  NAND4X0 U4304 ( .IN1(n5724), .IN2(n3805), .IN3(n3844), .IN4(n3803), .QN(
        n5045) );
  INVX0 U4305 ( .INP(n5073), .ZN(n5048) );
  INVX0 U4306 ( .INP(n5032), .ZN(n4427) );
  NAND2X0 U4307 ( .IN1(n5720), .IN2(n3844), .QN(n5032) );
  INVX0 U4308 ( .INP(n5039), .ZN(n5030) );
  NAND2X0 U4309 ( .IN1(n4420), .IN2(\r150/A[3] ), .QN(n5039) );
  INVX0 U4310 ( .INP(n4582), .ZN(n4420) );
  AO222X1 U4311 ( .IN1(n4519), .IN2(n5099), .IN3(n4523), .IN4(n5100), .IN5(
        n5101), .IN6(n4522), .Q(n5096) );
  AO222X1 U4312 ( .IN1(n4554), .IN2(n5102), .IN3(n4557), .IN4(n5103), .IN5(
        n5104), .IN6(n4556), .Q(n5100) );
  AO222X1 U4313 ( .IN1(n4583), .IN2(n5105), .IN3(n5106), .IN4(n4588), .IN5(
        n5107), .IN6(n4586), .Q(n5103) );
  AO222X1 U4314 ( .IN1(n4621), .IN2(n5108), .IN3(n4624), .IN4(n5109), .IN5(
        n5110), .IN6(n4591), .Q(n5106) );
  AO222X1 U4315 ( .IN1(n4654), .IN2(n5111), .IN3(n4658), .IN4(n5112), .IN5(
        n4656), .IN6(n5113), .Q(n5109) );
  AO222X1 U4316 ( .IN1(n4688), .IN2(n5114), .IN3(n4692), .IN4(n5115), .IN5(
        n5116), .IN6(n4691), .Q(n5112) );
  AO222X1 U4317 ( .IN1(n4724), .IN2(n5117), .IN3(n4727), .IN4(n5118), .IN5(
        n5119), .IN6(n4726), .Q(n5115) );
  AO222X1 U4318 ( .IN1(n4758), .IN2(n5120), .IN3(n4762), .IN4(n5121), .IN5(
        n5122), .IN6(n4761), .Q(n5118) );
  AO222X1 U4319 ( .IN1(n4797), .IN2(n5123), .IN3(n4753), .IN4(n5124), .IN5(
        n5125), .IN6(n4720), .Q(n5121) );
  AO222X1 U4320 ( .IN1(n4832), .IN2(n5126), .IN3(n4836), .IN4(n5127), .IN5(
        n4834), .IN6(n5128), .Q(n5124) );
  AO222X1 U4321 ( .IN1(n4876), .IN2(n5129), .IN3(n4880), .IN4(n5130), .IN5(
        n5131), .IN6(n4879), .Q(n5127) );
  AO222X1 U4322 ( .IN1(n4926), .IN2(n5132), .IN3(n4930), .IN4(n5133), .IN5(
        n4928), .IN6(n5134), .Q(n5130) );
  AO222X1 U4323 ( .IN1(n4970), .IN2(n5135), .IN3(n4974), .IN4(n5136), .IN5(
        n5137), .IN6(n4973), .Q(n5133) );
  AO22X1 U4324 ( .IN1(n4999), .IN2(n4265), .IN3(n5000), .IN4(n4266), .Q(n5136)
         );
  AND2X1 U4325 ( .IN1(n4489), .IN2(n4449), .Q(n4898) );
  AO222X1 U4326 ( .IN1(n5090), .IN2(n4488), .IN3(n4515), .IN4(n5138), .IN5(
        n4517), .IN6(n5091), .Q(n5095) );
  AO222X1 U4327 ( .IN1(n4549), .IN2(n5139), .IN3(n4551), .IN4(n5140), .IN5(
        n5141), .IN6(n4522), .Q(n5091) );
  AO222X1 U4328 ( .IN1(n5140), .IN2(n4522), .IN3(n4549), .IN4(n5142), .IN5(
        n4551), .IN6(n5139), .Q(n5138) );
  AO222X1 U4329 ( .IN1(n4589), .IN2(n5143), .IN3(n4592), .IN4(n5144), .IN5(
        n5145), .IN6(n4591), .Q(n5139) );
  AO222X1 U4330 ( .IN1(n5144), .IN2(n4591), .IN3(n4589), .IN4(n5146), .IN5(
        n4592), .IN6(n5143), .Q(n5142) );
  AO222X1 U4331 ( .IN1(n4557), .IN2(n5147), .IN3(n4619), .IN4(n5148), .IN5(
        n5149), .IN6(n4618), .Q(n5143) );
  AO222X1 U4332 ( .IN1(n5148), .IN2(n4618), .IN3(n4557), .IN4(n5150), .IN5(
        n4619), .IN6(n5147), .Q(n5146) );
  AO222X1 U4333 ( .IN1(n4649), .IN2(n5151), .IN3(n4652), .IN4(n5152), .IN5(
        n5153), .IN6(n4651), .Q(n5147) );
  AO222X1 U4334 ( .IN1(n5152), .IN2(n4651), .IN3(n4649), .IN4(n5154), .IN5(
        n4652), .IN6(n5151), .Q(n5150) );
  AO222X1 U4335 ( .IN1(n4683), .IN2(n5155), .IN3(n4686), .IN4(n5156), .IN5(
        n5157), .IN6(n4685), .Q(n5151) );
  AO222X1 U4336 ( .IN1(n4685), .IN2(n5156), .IN3(n5158), .IN4(n4683), .IN5(
        n5155), .IN6(n4686), .Q(n5154) );
  AO222X1 U4337 ( .IN1(n4718), .IN2(n5159), .IN3(n4721), .IN4(n5160), .IN5(
        n5161), .IN6(n4720), .Q(n5155) );
  AO221X1 U4338 ( .IN1(n5159), .IN2(n4721), .IN3(n4720), .IN4(n5160), .IN5(
        n5162), .Q(n5158) );
  OAI22X1 U4339 ( .IN1(n5163), .IN2(n5164), .IN3(n5165), .IN4(n4879), .QN(
        n5162) );
  AOI222X1 U4340 ( .IN1(n5166), .IN2(n4756), .IN3(n5167), .IN4(n4753), .IN5(
        n4755), .IN6(n5168), .QN(n5165) );
  AO22X1 U4341 ( .IN1(n5169), .IN2(n4789), .IN3(n5170), .IN4(n4792), .Q(n5167)
         );
  AO222X1 U4342 ( .IN1(n5171), .IN2(n4828), .IN3(n5172), .IN4(n4826), .IN5(
        n4761), .IN6(n5173), .Q(n5169) );
  AO222X1 U4343 ( .IN1(n5174), .IN2(n4869), .IN3(n5175), .IN4(n4866), .IN5(
        n5176), .IN6(n4868), .Q(n5172) );
  AO222X1 U4344 ( .IN1(n5177), .IN2(n4920), .IN3(n5178), .IN4(n4916), .IN5(
        n4919), .IN6(n5179), .Q(n5175) );
  AO222X1 U4345 ( .IN1(n5180), .IN2(n4966), .IN3(n5181), .IN4(n4727), .IN5(
        n4965), .IN6(n5182), .Q(n5178) );
  AO22X1 U4346 ( .IN1(n4327), .IN2(n5002), .IN3(n4325), .IN4(n5004), .Q(n5181)
         );
  NAND2X0 U4347 ( .IN1(n4876), .IN2(n5183), .QN(n5164) );
  AO222X1 U4348 ( .IN1(n4753), .IN2(n5166), .IN3(n4756), .IN4(n5168), .IN5(
        n5184), .IN6(n4755), .Q(n5159) );
  AO222X1 U4349 ( .IN1(n4789), .IN2(n5170), .IN3(n4792), .IN4(n5183), .IN5(
        n5185), .IN6(n4791), .Q(n5166) );
  AO222X1 U4350 ( .IN1(n4826), .IN2(n5171), .IN3(n4828), .IN4(n5173), .IN5(
        n5186), .IN6(n4761), .Q(n5170) );
  AO222X1 U4351 ( .IN1(n4866), .IN2(n5174), .IN3(n4869), .IN4(n5176), .IN5(
        n4868), .IN6(n5187), .Q(n5171) );
  AO222X1 U4352 ( .IN1(n4916), .IN2(n5177), .IN3(n4920), .IN4(n5179), .IN5(
        n5188), .IN6(n4919), .Q(n5174) );
  AO222X1 U4353 ( .IN1(n4727), .IN2(n5180), .IN3(n4966), .IN4(n5182), .IN5(
        n5189), .IN6(n4965), .Q(n5177) );
  AO222X1 U4354 ( .IN1(n5002), .IN2(n4328), .IN3(n5003), .IN4(n4325), .IN5(
        n5004), .IN6(n4327), .Q(n5180) );
  NOR2X0 U4355 ( .IN1(n5092), .IN2(n5017), .QN(n4447) );
  AO222X1 U4356 ( .IN1(n4517), .IN2(n5076), .IN3(n4516), .IN4(n4488), .IN5(
        n4515), .IN6(n5090), .Q(n4453) );
  AO222X1 U4357 ( .IN1(n4549), .IN2(n5140), .IN3(n5190), .IN4(n4522), .IN5(
        n4551), .IN6(n5141), .Q(n5090) );
  AO222X1 U4358 ( .IN1(n5191), .IN2(n4591), .IN3(n4589), .IN4(n5144), .IN5(
        n4592), .IN6(n5145), .Q(n5140) );
  AO222X1 U4359 ( .IN1(n5192), .IN2(n4618), .IN3(n4557), .IN4(n5148), .IN5(
        n4619), .IN6(n5149), .Q(n5144) );
  AO222X1 U4360 ( .IN1(n5193), .IN2(n4651), .IN3(n4649), .IN4(n5152), .IN5(
        n4652), .IN6(n5153), .Q(n5148) );
  AO222X1 U4361 ( .IN1(n5194), .IN2(n4685), .IN3(n4683), .IN4(n5156), .IN5(
        n4686), .IN6(n5157), .Q(n5152) );
  AO222X1 U4362 ( .IN1(n5195), .IN2(n4720), .IN3(n4718), .IN4(n5160), .IN5(
        n4721), .IN6(n5161), .Q(n5156) );
  AO222X1 U4363 ( .IN1(n5196), .IN2(n4755), .IN3(n4753), .IN4(n5168), .IN5(
        n4756), .IN6(n5184), .Q(n5160) );
  AO222X1 U4364 ( .IN1(n5197), .IN2(n4791), .IN3(n4789), .IN4(n5183), .IN5(
        n4792), .IN6(n5185), .Q(n5168) );
  AO222X1 U4365 ( .IN1(n5198), .IN2(n4761), .IN3(n4826), .IN4(n5173), .IN5(
        n4828), .IN6(n5186), .Q(n5183) );
  AO222X1 U4366 ( .IN1(n4868), .IN2(n5199), .IN3(n4866), .IN4(n5176), .IN5(
        n4869), .IN6(n5187), .Q(n5173) );
  AO222X1 U4367 ( .IN1(n5200), .IN2(n4919), .IN3(n4916), .IN4(n5179), .IN5(
        n4920), .IN6(n5188), .Q(n5176) );
  AO222X1 U4368 ( .IN1(n5201), .IN2(n4965), .IN3(n4727), .IN4(n5182), .IN5(
        n4966), .IN6(n5189), .Q(n5179) );
  AO222X1 U4369 ( .IN1(n5002), .IN2(n4329), .IN3(n5003), .IN4(n4327), .IN5(
        n5004), .IN6(n4328), .Q(n5182) );
  AO222X1 U4370 ( .IN1(n4551), .IN2(n5077), .IN3(n4550), .IN4(n4522), .IN5(
        n4549), .IN6(n5190), .Q(n4516) );
  AO222X1 U4371 ( .IN1(n4592), .IN2(n5078), .IN3(n4590), .IN4(n4591), .IN5(
        n4589), .IN6(n5202), .Q(n4550) );
  AO222X1 U4372 ( .IN1(n4619), .IN2(n5079), .IN3(n4617), .IN4(n4618), .IN5(
        n4557), .IN6(n5203), .Q(n4590) );
  AO222X1 U4373 ( .IN1(n4652), .IN2(n5080), .IN3(n4650), .IN4(n4651), .IN5(
        n4649), .IN6(n5204), .Q(n4617) );
  AO222X1 U4374 ( .IN1(n4686), .IN2(n5081), .IN3(n4684), .IN4(n4685), .IN5(
        n4683), .IN6(n5205), .Q(n4650) );
  AO222X1 U4375 ( .IN1(n4721), .IN2(n5082), .IN3(n4719), .IN4(n4720), .IN5(
        n4718), .IN6(n5206), .Q(n4684) );
  AO222X1 U4376 ( .IN1(n4756), .IN2(n5083), .IN3(n4754), .IN4(n4755), .IN5(
        n4753), .IN6(n5207), .Q(n4719) );
  AO222X1 U4377 ( .IN1(n4792), .IN2(n5084), .IN3(n4790), .IN4(n4791), .IN5(
        n4789), .IN6(n5208), .Q(n4754) );
  AO222X1 U4378 ( .IN1(n4828), .IN2(n5085), .IN3(n4827), .IN4(n4761), .IN5(
        n4826), .IN6(n5209), .Q(n4790) );
  AO222X1 U4379 ( .IN1(n4869), .IN2(n5086), .IN3(n4868), .IN4(n4867), .IN5(
        n4866), .IN6(n5210), .Q(n4827) );
  AO222X1 U4380 ( .IN1(n4920), .IN2(n5087), .IN3(n4917), .IN4(n4919), .IN5(
        n4916), .IN6(n5211), .Q(n4867) );
  AO222X1 U4381 ( .IN1(n4966), .IN2(n5088), .IN3(n4963), .IN4(n4965), .IN5(
        n4727), .IN6(n5212), .Q(n4917) );
  AO222X1 U4382 ( .IN1(n5002), .IN2(n4355), .IN3(n5003), .IN4(n4353), .IN5(
        n5004), .IN6(n4354), .Q(n4963) );
  AO222X1 U4383 ( .IN1(n4551), .IN2(n5190), .IN3(n5077), .IN4(n4522), .IN5(
        n4549), .IN6(n5141), .Q(n5076) );
  AO222X1 U4384 ( .IN1(n5213), .IN2(n4591), .IN3(n4592), .IN4(n5191), .IN5(
        n4589), .IN6(n5145), .Q(n5141) );
  AO222X1 U4385 ( .IN1(n5214), .IN2(n4618), .IN3(n4619), .IN4(n5192), .IN5(
        n4557), .IN6(n5149), .Q(n5145) );
  AO222X1 U4386 ( .IN1(n5215), .IN2(n4651), .IN3(n4652), .IN4(n5193), .IN5(
        n4649), .IN6(n5153), .Q(n5149) );
  AO222X1 U4387 ( .IN1(n4683), .IN2(n5157), .IN3(n4686), .IN4(n5194), .IN5(
        n5216), .IN6(n4685), .Q(n5153) );
  AO222X1 U4388 ( .IN1(n4718), .IN2(n5161), .IN3(n4721), .IN4(n5195), .IN5(
        n5217), .IN6(n4720), .Q(n5157) );
  AO222X1 U4389 ( .IN1(n4753), .IN2(n5184), .IN3(n4756), .IN4(n5196), .IN5(
        n4755), .IN6(n5218), .Q(n5161) );
  AO222X1 U4390 ( .IN1(n4789), .IN2(n5185), .IN3(n4792), .IN4(n5197), .IN5(
        n5219), .IN6(n4791), .Q(n5184) );
  AO222X1 U4391 ( .IN1(n4826), .IN2(n5186), .IN3(n4828), .IN4(n5198), .IN5(
        n5220), .IN6(n4761), .Q(n5185) );
  AO222X1 U4392 ( .IN1(n4866), .IN2(n5187), .IN3(n4869), .IN4(n5199), .IN5(
        n4868), .IN6(n5221), .Q(n5186) );
  AO222X1 U4393 ( .IN1(n4916), .IN2(n5188), .IN3(n4920), .IN4(n5200), .IN5(
        n5222), .IN6(n4919), .Q(n5187) );
  AO222X1 U4394 ( .IN1(n4727), .IN2(n5189), .IN3(n4966), .IN4(n5201), .IN5(
        n5223), .IN6(n4965), .Q(n5188) );
  AO222X1 U4395 ( .IN1(n5002), .IN2(n4330), .IN3(n5003), .IN4(n4328), .IN5(
        n5004), .IN6(n4329), .Q(n5189) );
  AO222X1 U4396 ( .IN1(n4592), .IN2(n5202), .IN3(n5078), .IN4(n4591), .IN5(
        n4589), .IN6(n5213), .Q(n5077) );
  AO222X1 U4397 ( .IN1(n4619), .IN2(n5203), .IN3(n5079), .IN4(n4618), .IN5(
        n4557), .IN6(n5224), .Q(n5078) );
  AO222X1 U4398 ( .IN1(n4652), .IN2(n5204), .IN3(n5080), .IN4(n4651), .IN5(
        n4649), .IN6(n5225), .Q(n5079) );
  AO222X1 U4399 ( .IN1(n4686), .IN2(n5205), .IN3(n5081), .IN4(n4685), .IN5(
        n4683), .IN6(n5226), .Q(n5080) );
  AO222X1 U4400 ( .IN1(n4721), .IN2(n5206), .IN3(n5082), .IN4(n4720), .IN5(
        n4718), .IN6(n5227), .Q(n5081) );
  AO222X1 U4401 ( .IN1(n4756), .IN2(n5207), .IN3(n5083), .IN4(n4755), .IN5(
        n4753), .IN6(n5228), .Q(n5082) );
  AO222X1 U4402 ( .IN1(n4792), .IN2(n5208), .IN3(n5084), .IN4(n4791), .IN5(
        n4789), .IN6(n5229), .Q(n5083) );
  AO222X1 U4403 ( .IN1(n4828), .IN2(n5209), .IN3(n5085), .IN4(n4761), .IN5(
        n4826), .IN6(n5230), .Q(n5084) );
  AO222X1 U4404 ( .IN1(n4869), .IN2(n5210), .IN3(n4868), .IN4(n5086), .IN5(
        n4866), .IN6(n5231), .Q(n5085) );
  AO222X1 U4405 ( .IN1(n4920), .IN2(n5211), .IN3(n5087), .IN4(n4919), .IN5(
        n4916), .IN6(n5232), .Q(n5086) );
  AO222X1 U4406 ( .IN1(n4966), .IN2(n5212), .IN3(n5088), .IN4(n4965), .IN5(
        n4727), .IN6(n5233), .Q(n5087) );
  AO222X1 U4407 ( .IN1(n5002), .IN2(n4354), .IN3(n5003), .IN4(n4352), .IN5(
        n5004), .IN6(n4353), .Q(n5088) );
  AO222X1 U4408 ( .IN1(n4589), .IN2(n5191), .IN3(n5202), .IN4(n4591), .IN5(
        n4592), .IN6(n5213), .Q(n5190) );
  AO222X1 U4409 ( .IN1(n5224), .IN2(n4618), .IN3(n4619), .IN4(n5234), .IN5(
        n4557), .IN6(n5214), .Q(n5213) );
  NOR2X0 U4410 ( .IN1(n4591), .IN2(n4589), .QN(n4592) );
  AO222X1 U4411 ( .IN1(n4557), .IN2(n5234), .IN3(n5203), .IN4(n4618), .IN5(
        n4619), .IN6(n5224), .Q(n5202) );
  AO222X1 U4412 ( .IN1(n5225), .IN2(n4651), .IN3(n4652), .IN4(n5235), .IN5(
        n4649), .IN6(n5236), .Q(n5224) );
  AO222X1 U4413 ( .IN1(n4649), .IN2(n5235), .IN3(n5204), .IN4(n4651), .IN5(
        n4652), .IN6(n5225), .Q(n5203) );
  AO222X1 U4414 ( .IN1(n5226), .IN2(n4685), .IN3(n4686), .IN4(n5237), .IN5(
        n4683), .IN6(n5238), .Q(n5225) );
  AO222X1 U4415 ( .IN1(n4683), .IN2(n5237), .IN3(n5205), .IN4(n4685), .IN5(
        n4686), .IN6(n5226), .Q(n5204) );
  AO222X1 U4416 ( .IN1(n5227), .IN2(n4720), .IN3(n4721), .IN4(n5239), .IN5(
        n4718), .IN6(n5240), .Q(n5226) );
  AO222X1 U4417 ( .IN1(n4718), .IN2(n5239), .IN3(n5206), .IN4(n4720), .IN5(
        n4721), .IN6(n5227), .Q(n5205) );
  AO222X1 U4418 ( .IN1(n5228), .IN2(n4755), .IN3(n4756), .IN4(n5241), .IN5(
        n4753), .IN6(n5242), .Q(n5227) );
  AO222X1 U4419 ( .IN1(n4753), .IN2(n5241), .IN3(n5207), .IN4(n4755), .IN5(
        n4756), .IN6(n5228), .Q(n5206) );
  AO222X1 U4420 ( .IN1(n5229), .IN2(n4791), .IN3(n4792), .IN4(n5243), .IN5(
        n4789), .IN6(n5244), .Q(n5228) );
  AO222X1 U4421 ( .IN1(n4789), .IN2(n5243), .IN3(n5208), .IN4(n4791), .IN5(
        n4792), .IN6(n5229), .Q(n5207) );
  AO222X1 U4422 ( .IN1(n5230), .IN2(n4761), .IN3(n4828), .IN4(n5245), .IN5(
        n4826), .IN6(n5246), .Q(n5229) );
  AO222X1 U4423 ( .IN1(n4826), .IN2(n5245), .IN3(n5209), .IN4(n4761), .IN5(
        n4828), .IN6(n5230), .Q(n5208) );
  AO222X1 U4424 ( .IN1(n4868), .IN2(n5231), .IN3(n4869), .IN4(n5247), .IN5(
        n4866), .IN6(n5248), .Q(n5230) );
  AO222X1 U4425 ( .IN1(n4866), .IN2(n5247), .IN3(n4868), .IN4(n5210), .IN5(
        n4869), .IN6(n5231), .Q(n5209) );
  AO222X1 U4426 ( .IN1(n5232), .IN2(n4919), .IN3(n4920), .IN4(n5249), .IN5(
        n4916), .IN6(n5250), .Q(n5231) );
  AO222X1 U4427 ( .IN1(n4916), .IN2(n5249), .IN3(n5211), .IN4(n4919), .IN5(
        n4920), .IN6(n5232), .Q(n5210) );
  AO222X1 U4428 ( .IN1(n5233), .IN2(n4965), .IN3(n4966), .IN4(n5251), .IN5(
        n4727), .IN6(n5252), .Q(n5232) );
  AO222X1 U4429 ( .IN1(n4727), .IN2(n5251), .IN3(n5212), .IN4(n4965), .IN5(
        n4966), .IN6(n5233), .Q(n5211) );
  AO222X1 U4430 ( .IN1(n5002), .IN2(n4352), .IN3(n5003), .IN4(n4350), .IN5(
        n5004), .IN6(n4351), .Q(n5233) );
  AO222X1 U4431 ( .IN1(n5002), .IN2(n4353), .IN3(n5003), .IN4(n4351), .IN5(
        n5004), .IN6(n4352), .Q(n5212) );
  AO222X1 U4432 ( .IN1(n4557), .IN2(n5192), .IN3(n5234), .IN4(n4618), .IN5(
        n4619), .IN6(n5214), .Q(n5191) );
  AO222X1 U4433 ( .IN1(n5236), .IN2(n4651), .IN3(n4652), .IN4(n5253), .IN5(
        n4649), .IN6(n5215), .Q(n5214) );
  NOR2X0 U4434 ( .IN1(n4557), .IN2(n4618), .QN(n4619) );
  AO222X1 U4435 ( .IN1(n4649), .IN2(n5253), .IN3(n5235), .IN4(n4651), .IN5(
        n4652), .IN6(n5236), .Q(n5234) );
  AO222X1 U4436 ( .IN1(n5238), .IN2(n4685), .IN3(n4686), .IN4(n5254), .IN5(
        n4683), .IN6(n5255), .Q(n5236) );
  AO222X1 U4437 ( .IN1(n4683), .IN2(n5254), .IN3(n5237), .IN4(n4685), .IN5(
        n4686), .IN6(n5238), .Q(n5235) );
  AO222X1 U4438 ( .IN1(n5240), .IN2(n4720), .IN3(n4721), .IN4(n5256), .IN5(
        n4718), .IN6(n5257), .Q(n5238) );
  AO222X1 U4439 ( .IN1(n4718), .IN2(n5256), .IN3(n5239), .IN4(n4720), .IN5(
        n4721), .IN6(n5240), .Q(n5237) );
  AO222X1 U4440 ( .IN1(n5242), .IN2(n4755), .IN3(n4756), .IN4(n5258), .IN5(
        n4753), .IN6(n5259), .Q(n5240) );
  AO222X1 U4441 ( .IN1(n4753), .IN2(n5258), .IN3(n5241), .IN4(n4755), .IN5(
        n4756), .IN6(n5242), .Q(n5239) );
  AO222X1 U4442 ( .IN1(n5244), .IN2(n4791), .IN3(n4792), .IN4(n5260), .IN5(
        n4789), .IN6(n5261), .Q(n5242) );
  AO222X1 U4443 ( .IN1(n4789), .IN2(n5260), .IN3(n5243), .IN4(n4791), .IN5(
        n4792), .IN6(n5244), .Q(n5241) );
  AO222X1 U4444 ( .IN1(n5246), .IN2(n4761), .IN3(n4828), .IN4(n5262), .IN5(
        n4826), .IN6(n5263), .Q(n5244) );
  AO222X1 U4445 ( .IN1(n4826), .IN2(n5262), .IN3(n5245), .IN4(n4761), .IN5(
        n4828), .IN6(n5246), .Q(n5243) );
  AO222X1 U4446 ( .IN1(n4868), .IN2(n5248), .IN3(n4869), .IN4(n5264), .IN5(
        n4866), .IN6(n5265), .Q(n5246) );
  AO222X1 U4447 ( .IN1(n4866), .IN2(n5264), .IN3(n4868), .IN4(n5247), .IN5(
        n4869), .IN6(n5248), .Q(n5245) );
  AO222X1 U4448 ( .IN1(n5250), .IN2(n4919), .IN3(n4920), .IN4(n5266), .IN5(
        n4916), .IN6(n5267), .Q(n5248) );
  AO222X1 U4449 ( .IN1(n4916), .IN2(n5266), .IN3(n5249), .IN4(n4919), .IN5(
        n4920), .IN6(n5250), .Q(n5247) );
  AO222X1 U4450 ( .IN1(n5252), .IN2(n4965), .IN3(n4966), .IN4(n5268), .IN5(
        n4727), .IN6(n5269), .Q(n5250) );
  AO222X1 U4451 ( .IN1(n4727), .IN2(n5268), .IN3(n5251), .IN4(n4965), .IN5(
        n4966), .IN6(n5252), .Q(n5249) );
  AO222X1 U4452 ( .IN1(n5002), .IN2(n4350), .IN3(n5003), .IN4(n4348), .IN5(
        n5004), .IN6(n4349), .Q(n5252) );
  AO222X1 U4453 ( .IN1(n5002), .IN2(n4351), .IN3(n5003), .IN4(n4349), .IN5(
        n5004), .IN6(n4350), .Q(n5251) );
  AO222X1 U4454 ( .IN1(n4649), .IN2(n5193), .IN3(n5253), .IN4(n4651), .IN5(
        n4652), .IN6(n5215), .Q(n5192) );
  AO222X1 U4455 ( .IN1(n5255), .IN2(n4685), .IN3(n4686), .IN4(n5270), .IN5(
        n4683), .IN6(n5216), .Q(n5215) );
  NOR2X0 U4456 ( .IN1(n4651), .IN2(n4649), .QN(n4652) );
  AO222X1 U4457 ( .IN1(n4683), .IN2(n5270), .IN3(n5254), .IN4(n4685), .IN5(
        n4686), .IN6(n5255), .Q(n5253) );
  AO222X1 U4458 ( .IN1(n5257), .IN2(n4720), .IN3(n4721), .IN4(n5271), .IN5(
        n4718), .IN6(n5272), .Q(n5255) );
  AO222X1 U4459 ( .IN1(n4718), .IN2(n5271), .IN3(n5256), .IN4(n4720), .IN5(
        n4721), .IN6(n5257), .Q(n5254) );
  AO222X1 U4460 ( .IN1(n5259), .IN2(n4755), .IN3(n4756), .IN4(n5273), .IN5(
        n4753), .IN6(n5274), .Q(n5257) );
  AO222X1 U4461 ( .IN1(n4753), .IN2(n5273), .IN3(n5258), .IN4(n4755), .IN5(
        n4756), .IN6(n5259), .Q(n5256) );
  AO222X1 U4462 ( .IN1(n5261), .IN2(n4791), .IN3(n4792), .IN4(n5275), .IN5(
        n4789), .IN6(n5276), .Q(n5259) );
  AO222X1 U4463 ( .IN1(n4789), .IN2(n5275), .IN3(n5260), .IN4(n4791), .IN5(
        n4792), .IN6(n5261), .Q(n5258) );
  AO222X1 U4464 ( .IN1(n5263), .IN2(n4761), .IN3(n4828), .IN4(n5277), .IN5(
        n4826), .IN6(n5278), .Q(n5261) );
  AO222X1 U4465 ( .IN1(n4826), .IN2(n5277), .IN3(n5262), .IN4(n4761), .IN5(
        n4828), .IN6(n5263), .Q(n5260) );
  AO222X1 U4466 ( .IN1(n4868), .IN2(n5265), .IN3(n4869), .IN4(n5279), .IN5(
        n4866), .IN6(n5280), .Q(n5263) );
  AO222X1 U4467 ( .IN1(n4866), .IN2(n5279), .IN3(n4868), .IN4(n5264), .IN5(
        n4869), .IN6(n5265), .Q(n5262) );
  AO222X1 U4468 ( .IN1(n5267), .IN2(n4919), .IN3(n4920), .IN4(n5281), .IN5(
        n4916), .IN6(n5282), .Q(n5265) );
  AO222X1 U4469 ( .IN1(n4916), .IN2(n5281), .IN3(n5266), .IN4(n4919), .IN5(
        n4920), .IN6(n5267), .Q(n5264) );
  AO222X1 U4470 ( .IN1(n5269), .IN2(n4965), .IN3(n4966), .IN4(n5283), .IN5(
        n4727), .IN6(n5284), .Q(n5267) );
  AO222X1 U4471 ( .IN1(n4727), .IN2(n5283), .IN3(n5268), .IN4(n4965), .IN5(
        n4966), .IN6(n5269), .Q(n5266) );
  AO222X1 U4472 ( .IN1(n5002), .IN2(n4348), .IN3(n5003), .IN4(n4346), .IN5(
        n5004), .IN6(n4347), .Q(n5269) );
  AO222X1 U4473 ( .IN1(n5002), .IN2(n4349), .IN3(n5003), .IN4(n4347), .IN5(
        n5004), .IN6(n4348), .Q(n5268) );
  AO222X1 U4474 ( .IN1(n4683), .IN2(n5194), .IN3(n5270), .IN4(n4685), .IN5(
        n4686), .IN6(n5216), .Q(n5193) );
  AO222X1 U4475 ( .IN1(n5272), .IN2(n4720), .IN3(n4721), .IN4(n5285), .IN5(
        n4718), .IN6(n5217), .Q(n5216) );
  NOR2X0 U4476 ( .IN1(n4685), .IN2(n4683), .QN(n4686) );
  AO222X1 U4477 ( .IN1(n4718), .IN2(n5285), .IN3(n5271), .IN4(n4720), .IN5(
        n4721), .IN6(n5272), .Q(n5270) );
  AO222X1 U4478 ( .IN1(n5274), .IN2(n4755), .IN3(n4756), .IN4(n5286), .IN5(
        n4753), .IN6(n5287), .Q(n5272) );
  AO222X1 U4479 ( .IN1(n4753), .IN2(n5286), .IN3(n5273), .IN4(n4755), .IN5(
        n4756), .IN6(n5274), .Q(n5271) );
  AO222X1 U4480 ( .IN1(n5276), .IN2(n4791), .IN3(n4792), .IN4(n5288), .IN5(
        n4789), .IN6(n5289), .Q(n5274) );
  AO222X1 U4481 ( .IN1(n4789), .IN2(n5288), .IN3(n5275), .IN4(n4791), .IN5(
        n4792), .IN6(n5276), .Q(n5273) );
  AO222X1 U4482 ( .IN1(n5278), .IN2(n4761), .IN3(n4828), .IN4(n5290), .IN5(
        n4826), .IN6(n5291), .Q(n5276) );
  AO222X1 U4483 ( .IN1(n4826), .IN2(n5290), .IN3(n5277), .IN4(n4761), .IN5(
        n4828), .IN6(n5278), .Q(n5275) );
  AO222X1 U4484 ( .IN1(n4868), .IN2(n5280), .IN3(n4869), .IN4(n5292), .IN5(
        n4866), .IN6(n5293), .Q(n5278) );
  AO222X1 U4485 ( .IN1(n4866), .IN2(n5292), .IN3(n4868), .IN4(n5279), .IN5(
        n4869), .IN6(n5280), .Q(n5277) );
  AO222X1 U4486 ( .IN1(n5282), .IN2(n4919), .IN3(n4920), .IN4(n5294), .IN5(
        n4916), .IN6(n5295), .Q(n5280) );
  AO222X1 U4487 ( .IN1(n4916), .IN2(n5294), .IN3(n5281), .IN4(n4919), .IN5(
        n4920), .IN6(n5282), .Q(n5279) );
  AO222X1 U4488 ( .IN1(n5284), .IN2(n4965), .IN3(n4966), .IN4(n5296), .IN5(
        n4727), .IN6(n5297), .Q(n5282) );
  AO222X1 U4489 ( .IN1(n4727), .IN2(n5296), .IN3(n5283), .IN4(n4965), .IN5(
        n4966), .IN6(n5284), .Q(n5281) );
  AO222X1 U4490 ( .IN1(n5002), .IN2(n4346), .IN3(n5003), .IN4(n4344), .IN5(
        n5004), .IN6(n4345), .Q(n5284) );
  AO222X1 U4491 ( .IN1(n5002), .IN2(n4347), .IN3(n5003), .IN4(n4345), .IN5(
        n5004), .IN6(n4346), .Q(n5283) );
  AO222X1 U4492 ( .IN1(n5285), .IN2(n4720), .IN3(n4718), .IN4(n5195), .IN5(
        n4721), .IN6(n5217), .Q(n5194) );
  AO222X1 U4493 ( .IN1(n4755), .IN2(n5287), .IN3(n4756), .IN4(n5298), .IN5(
        n4753), .IN6(n5218), .Q(n5217) );
  NOR2X0 U4494 ( .IN1(n4720), .IN2(n4718), .QN(n4721) );
  AO222X1 U4495 ( .IN1(n5298), .IN2(n4755), .IN3(n4753), .IN4(n5196), .IN5(
        n4756), .IN6(n5218), .Q(n5195) );
  AO222X1 U4496 ( .IN1(n5299), .IN2(n4791), .IN3(n4792), .IN4(n5300), .IN5(
        n4789), .IN6(n5219), .Q(n5218) );
  AO222X1 U4497 ( .IN1(n5300), .IN2(n4791), .IN3(n4789), .IN4(n5197), .IN5(
        n4792), .IN6(n5219), .Q(n5196) );
  AO222X1 U4498 ( .IN1(n5301), .IN2(n4761), .IN3(n4828), .IN4(n5302), .IN5(
        n4826), .IN6(n5220), .Q(n5219) );
  AO222X1 U4499 ( .IN1(n5302), .IN2(n4761), .IN3(n4826), .IN4(n5198), .IN5(
        n4828), .IN6(n5220), .Q(n5197) );
  AO222X1 U4500 ( .IN1(n4866), .IN2(n5221), .IN3(n4869), .IN4(n5303), .IN5(
        n4868), .IN6(n5304), .Q(n5220) );
  AO222X1 U4501 ( .IN1(n4868), .IN2(n5303), .IN3(n4866), .IN4(n5199), .IN5(
        n4869), .IN6(n5221), .Q(n5198) );
  AO222X1 U4502 ( .IN1(n4916), .IN2(n5222), .IN3(n4920), .IN4(n5305), .IN5(
        n5306), .IN6(n4919), .Q(n5221) );
  AO222X1 U4503 ( .IN1(n5305), .IN2(n4919), .IN3(n4916), .IN4(n5200), .IN5(
        n4920), .IN6(n5222), .Q(n5199) );
  AO222X1 U4504 ( .IN1(n4727), .IN2(n5223), .IN3(n4966), .IN4(n5307), .IN5(
        n5308), .IN6(n4965), .Q(n5222) );
  AO222X1 U4505 ( .IN1(n5307), .IN2(n4965), .IN3(n4727), .IN4(n5201), .IN5(
        n4966), .IN6(n5223), .Q(n5200) );
  AO222X1 U4506 ( .IN1(n5002), .IN2(n4332), .IN3(n5003), .IN4(n4330), .IN5(
        n5004), .IN6(n4331), .Q(n5223) );
  AO222X1 U4507 ( .IN1(n5002), .IN2(n4331), .IN3(n5003), .IN4(n4329), .IN5(
        n5004), .IN6(n4330), .Q(n5201) );
  INVX0 U4508 ( .INP(n4879), .ZN(n4718) );
  AO222X1 U4509 ( .IN1(n4753), .IN2(n5298), .IN3(n5286), .IN4(n4755), .IN5(
        n4756), .IN6(n5287), .Q(n5285) );
  AO222X1 U4510 ( .IN1(n5289), .IN2(n4791), .IN3(n4792), .IN4(n5309), .IN5(
        n4789), .IN6(n5299), .Q(n5287) );
  NOR2X0 U4511 ( .IN1(n4755), .IN2(n4753), .QN(n4756) );
  NAND3X0 U4512 ( .IN1(n5310), .IN2(n5311), .IN3(n5312), .QN(n4755) );
  OR2X1 U4513 ( .IN1(n5313), .IN2(n5314), .Q(n5312) );
  AO222X1 U4514 ( .IN1(n4789), .IN2(n5309), .IN3(n5288), .IN4(n4791), .IN5(
        n4792), .IN6(n5289), .Q(n5286) );
  AO222X1 U4515 ( .IN1(n5291), .IN2(n4761), .IN3(n4828), .IN4(n5315), .IN5(
        n4826), .IN6(n5316), .Q(n5289) );
  AO222X1 U4516 ( .IN1(n4826), .IN2(n5315), .IN3(n5290), .IN4(n4761), .IN5(
        n4828), .IN6(n5291), .Q(n5288) );
  AO222X1 U4517 ( .IN1(n4868), .IN2(n5293), .IN3(n4869), .IN4(n5317), .IN5(
        n4866), .IN6(n5318), .Q(n5291) );
  AO222X1 U4518 ( .IN1(n4866), .IN2(n5317), .IN3(n4868), .IN4(n5292), .IN5(
        n4869), .IN6(n5293), .Q(n5290) );
  AO222X1 U4519 ( .IN1(n5295), .IN2(n4919), .IN3(n4920), .IN4(n5319), .IN5(
        n4916), .IN6(n5320), .Q(n5293) );
  AO222X1 U4520 ( .IN1(n4916), .IN2(n5319), .IN3(n5294), .IN4(n4919), .IN5(
        n4920), .IN6(n5295), .Q(n5292) );
  AO222X1 U4521 ( .IN1(n5297), .IN2(n4965), .IN3(n4966), .IN4(n5321), .IN5(
        n4727), .IN6(n5322), .Q(n5295) );
  AO222X1 U4522 ( .IN1(n4727), .IN2(n5321), .IN3(n5296), .IN4(n4965), .IN5(
        n4966), .IN6(n5297), .Q(n5294) );
  AO222X1 U4523 ( .IN1(n5002), .IN2(n4344), .IN3(n5003), .IN4(n4342), .IN5(
        n5004), .IN6(n4343), .Q(n5297) );
  AO222X1 U4524 ( .IN1(n5002), .IN2(n4345), .IN3(n5003), .IN4(n4343), .IN5(
        n5004), .IN6(n4344), .Q(n5296) );
  AO222X1 U4525 ( .IN1(n4789), .IN2(n5300), .IN3(n5309), .IN4(n4791), .IN5(
        n4792), .IN6(n5299), .Q(n5298) );
  AO222X1 U4526 ( .IN1(n5316), .IN2(n4761), .IN3(n4828), .IN4(n5323), .IN5(
        n4826), .IN6(n5301), .Q(n5299) );
  NOR2X0 U4527 ( .IN1(n4791), .IN2(n4789), .QN(n4792) );
  INVX0 U4528 ( .INP(n4880), .ZN(n4791) );
  AO222X1 U4529 ( .IN1(n4826), .IN2(n5323), .IN3(n5315), .IN4(n4761), .IN5(
        n4828), .IN6(n5316), .Q(n5309) );
  AO222X1 U4530 ( .IN1(n4868), .IN2(n5318), .IN3(n4869), .IN4(n5324), .IN5(
        n4866), .IN6(n5325), .Q(n5316) );
  AO222X1 U4531 ( .IN1(n4866), .IN2(n5324), .IN3(n4868), .IN4(n5317), .IN5(
        n4869), .IN6(n5318), .Q(n5315) );
  AO222X1 U4532 ( .IN1(n5320), .IN2(n4919), .IN3(n4920), .IN4(n5326), .IN5(
        n4916), .IN6(n5327), .Q(n5318) );
  AO222X1 U4533 ( .IN1(n4916), .IN2(n5326), .IN3(n5319), .IN4(n4919), .IN5(
        n4920), .IN6(n5320), .Q(n5317) );
  AO222X1 U4534 ( .IN1(n5322), .IN2(n4965), .IN3(n4966), .IN4(n5328), .IN5(
        n4727), .IN6(n5329), .Q(n5320) );
  AO222X1 U4535 ( .IN1(n4727), .IN2(n5328), .IN3(n5321), .IN4(n4965), .IN5(
        n4966), .IN6(n5322), .Q(n5319) );
  AO222X1 U4536 ( .IN1(n5002), .IN2(n4342), .IN3(n5003), .IN4(n4340), .IN5(
        n5004), .IN6(n4341), .Q(n5322) );
  AO222X1 U4537 ( .IN1(n5002), .IN2(n4343), .IN3(n5003), .IN4(n4341), .IN5(
        n5004), .IN6(n4342), .Q(n5321) );
  AO222X1 U4538 ( .IN1(n4826), .IN2(n5302), .IN3(n5323), .IN4(n4761), .IN5(
        n4828), .IN6(n5301), .Q(n5300) );
  AO222X1 U4539 ( .IN1(n4868), .IN2(n5325), .IN3(n4869), .IN4(n5330), .IN5(
        n4866), .IN6(n5304), .Q(n5301) );
  NOR2X0 U4540 ( .IN1(n4761), .IN2(n4826), .QN(n4828) );
  AO222X1 U4541 ( .IN1(n4866), .IN2(n5330), .IN3(n4868), .IN4(n5324), .IN5(
        n4869), .IN6(n5325), .Q(n5323) );
  AO222X1 U4542 ( .IN1(n5327), .IN2(n4919), .IN3(n4920), .IN4(n5331), .IN5(
        n4916), .IN6(n5332), .Q(n5325) );
  AO222X1 U4543 ( .IN1(n4916), .IN2(n5331), .IN3(n5326), .IN4(n4919), .IN5(
        n4920), .IN6(n5327), .Q(n5324) );
  AO222X1 U4544 ( .IN1(n5329), .IN2(n4965), .IN3(n4966), .IN4(n5333), .IN5(
        n4727), .IN6(n5334), .Q(n5327) );
  AO222X1 U4545 ( .IN1(n4727), .IN2(n5333), .IN3(n5328), .IN4(n4965), .IN5(
        n4966), .IN6(n5329), .Q(n5326) );
  AO222X1 U4546 ( .IN1(n5002), .IN2(n4340), .IN3(n5003), .IN4(n4338), .IN5(
        n5004), .IN6(n4339), .Q(n5329) );
  AO222X1 U4547 ( .IN1(n5002), .IN2(n4341), .IN3(n5003), .IN4(n4339), .IN5(
        n5004), .IN6(n4340), .Q(n5328) );
  AO222X1 U4548 ( .IN1(n4866), .IN2(n5303), .IN3(n4868), .IN4(n5330), .IN5(
        n4869), .IN6(n5304), .Q(n5302) );
  AO222X1 U4549 ( .IN1(n5332), .IN2(n4919), .IN3(n4920), .IN4(n5335), .IN5(
        n4916), .IN6(n5306), .Q(n5304) );
  NOR2X0 U4550 ( .IN1(n5336), .IN2(n5337), .QN(n4869) );
  AO222X1 U4551 ( .IN1(n4916), .IN2(n5335), .IN3(n5331), .IN4(n4919), .IN5(
        n4920), .IN6(n5332), .Q(n5330) );
  AO222X1 U4552 ( .IN1(n5334), .IN2(n4965), .IN3(n4966), .IN4(n5338), .IN5(
        n4727), .IN6(n5339), .Q(n5332) );
  AO222X1 U4553 ( .IN1(n4727), .IN2(n5338), .IN3(n5333), .IN4(n4965), .IN5(
        n4966), .IN6(n5334), .Q(n5331) );
  AO222X1 U4554 ( .IN1(n5002), .IN2(n4338), .IN3(n5003), .IN4(n4336), .IN5(
        n5004), .IN6(n4337), .Q(n5334) );
  AO222X1 U4555 ( .IN1(n5002), .IN2(n4339), .IN3(n5003), .IN4(n4337), .IN5(
        n5004), .IN6(n4338), .Q(n5333) );
  NOR2X0 U4556 ( .IN1(n5337), .IN2(n4974), .QN(n4868) );
  AO222X1 U4557 ( .IN1(n5335), .IN2(n4919), .IN3(n4916), .IN4(n5305), .IN5(
        n4920), .IN6(n5306), .Q(n5303) );
  AO222X1 U4558 ( .IN1(n5339), .IN2(n4965), .IN3(n4966), .IN4(n5340), .IN5(
        n4727), .IN6(n5308), .Q(n5306) );
  NOR2X0 U4559 ( .IN1(n4919), .IN2(n4916), .QN(n4920) );
  AO222X1 U4560 ( .IN1(n5340), .IN2(n4965), .IN3(n4727), .IN4(n5307), .IN5(
        n4966), .IN6(n5308), .Q(n5305) );
  AO222X1 U4561 ( .IN1(n5002), .IN2(n4334), .IN3(n5003), .IN4(n4332), .IN5(
        n5004), .IN6(n4333), .Q(n5308) );
  AO222X1 U4562 ( .IN1(n5002), .IN2(n4333), .IN3(n5003), .IN4(n4331), .IN5(
        n5004), .IN6(n4332), .Q(n5307) );
  AO222X1 U4563 ( .IN1(n4727), .IN2(n5340), .IN3(n5338), .IN4(n4965), .IN5(
        n4966), .IN6(n5339), .Q(n5335) );
  AO222X1 U4564 ( .IN1(n5002), .IN2(n4336), .IN3(n5003), .IN4(n4334), .IN5(
        n5004), .IN6(n4335), .Q(n5339) );
  NOR2X0 U4565 ( .IN1(n4965), .IN2(n4727), .QN(n4966) );
  AO222X1 U4566 ( .IN1(n5002), .IN2(n4337), .IN3(n5003), .IN4(n4335), .IN5(
        n5004), .IN6(n4336), .Q(n5338) );
  AO222X1 U4567 ( .IN1(n5002), .IN2(n4335), .IN3(n5003), .IN4(n4333), .IN5(
        n5004), .IN6(n4334), .Q(n5340) );
  XOR2X1 U4568 ( .IN1(n5341), .IN2(n5342), .Q(n5004) );
  NOR2X0 U4569 ( .IN1(n5342), .IN2(n5341), .QN(n5003) );
  NOR2X0 U4570 ( .IN1(n5001), .IN2(n4692), .QN(n5002) );
  NOR2X0 U4571 ( .IN1(n5336), .IN2(n4586), .QN(n4866) );
  INVX0 U4572 ( .INP(n4973), .ZN(n4683) );
  INVX0 U4573 ( .INP(n4691), .ZN(n4589) );
  NOR2X0 U4574 ( .IN1(n4549), .IN2(n4522), .QN(n4551) );
  NOR2X0 U4575 ( .IN1(n4488), .IN2(n4515), .QN(n4517) );
  AND2X1 U4576 ( .IN1(n4942), .IN2(n4726), .Q(n4454) );
  INVX0 U4577 ( .INP(n5092), .ZN(n4942) );
  NAND2X0 U4578 ( .IN1(n5027), .IN2(n5343), .QN(n5092) );
  NOR4X0 U4579 ( .IN1(n5344), .IN2(n5075), .IN3(n3804), .IN4(n3843), .QN(n5027) );
  AND2X1 U4580 ( .IN1(n4485), .IN2(n4449), .Q(n4894) );
  AND2X1 U4581 ( .IN1(n5345), .IN2(n5343), .Q(n4449) );
  AO221X1 U4582 ( .IN1(N3826), .IN2(n4466), .IN3(n4459), .IN4(n4450), .IN5(
        n5346), .Q(n5062) );
  AO21X1 U4583 ( .IN1(N3720), .IN2(n4468), .IN3(n4469), .Q(n5346) );
  AO21X1 U4584 ( .IN1(n5347), .IN2(n4417), .IN3(n5033), .Q(n4469) );
  AND4X1 U4585 ( .IN1(n5348), .IN2(n5722), .IN3(n5349), .IN4(n5724), .Q(n5033)
         );
  AND2X1 U4586 ( .IN1(n4357), .IN2(n5344), .Q(n5349) );
  INVX0 U4587 ( .INP(n5014), .ZN(n5347) );
  NAND3X0 U4588 ( .IN1(n5723), .IN2(n4296), .IN3(n5350), .QN(n5014) );
  INVX0 U4589 ( .INP(n5725), .ZN(n4296) );
  AND3X1 U4590 ( .IN1(n3843), .IN2(n3804), .IN3(n5350), .Q(n4468) );
  AO222X1 U4591 ( .IN1(n4489), .IN2(n5093), .IN3(n4486), .IN4(n4488), .IN5(
        n4485), .IN6(n4490), .Q(n4450) );
  AO222X1 U4592 ( .IN1(n4523), .IN2(n5101), .IN3(n4524), .IN4(n4522), .IN5(
        n4519), .IN6(n5351), .Q(n4490) );
  NOR2X0 U4593 ( .IN1(n4488), .IN2(n4489), .QN(n4485) );
  OAI21X1 U4594 ( .IN1(n5352), .IN2(n5353), .IN3(n5354), .QN(n4488) );
  AO222X1 U4595 ( .IN1(n4519), .IN2(n4524), .IN3(n4520), .IN4(n4522), .IN5(
        n4523), .IN6(n5351), .Q(n4486) );
  AO222X1 U4596 ( .IN1(n4554), .IN2(n4558), .IN3(n4555), .IN4(n4556), .IN5(
        n4557), .IN6(n5355), .Q(n4520) );
  AO222X1 U4597 ( .IN1(n4583), .IN2(n4587), .IN3(n4584), .IN4(n4586), .IN5(
        n5356), .IN6(n4588), .Q(n4555) );
  AO222X1 U4598 ( .IN1(n4621), .IN2(n4625), .IN3(n4622), .IN4(n4591), .IN5(
        n4624), .IN6(n5357), .Q(n4584) );
  AO222X1 U4599 ( .IN1(n4654), .IN2(n4659), .IN3(n4656), .IN4(n4655), .IN5(
        n4658), .IN6(n5358), .Q(n4622) );
  AO222X1 U4600 ( .IN1(n4688), .IN2(n4693), .IN3(n4689), .IN4(n4691), .IN5(
        n4692), .IN6(n5359), .Q(n4655) );
  AO222X1 U4601 ( .IN1(n4724), .IN2(n4728), .IN3(n4725), .IN4(n4726), .IN5(
        n4727), .IN6(n5360), .Q(n4689) );
  AO222X1 U4602 ( .IN1(n4758), .IN2(n4763), .IN3(n4759), .IN4(n4761), .IN5(
        n4762), .IN6(n5361), .Q(n4725) );
  AO222X1 U4603 ( .IN1(n4797), .IN2(n4800), .IN3(n4798), .IN4(n4720), .IN5(
        n4753), .IN6(n5362), .Q(n4759) );
  AO222X1 U4604 ( .IN1(n4832), .IN2(n4837), .IN3(n4834), .IN4(n4833), .IN5(
        n4836), .IN6(n5363), .Q(n4798) );
  AO222X1 U4605 ( .IN1(n4876), .IN2(n4881), .IN3(n4877), .IN4(n4879), .IN5(
        n4880), .IN6(n5364), .Q(n4833) );
  AO222X1 U4606 ( .IN1(n4926), .IN2(n4931), .IN3(n4928), .IN4(n4927), .IN5(
        n4930), .IN6(n5365), .Q(n4877) );
  AO222X1 U4607 ( .IN1(n4970), .IN2(n4975), .IN3(n4971), .IN4(n4973), .IN5(
        n4974), .IN6(n5366), .Q(n4927) );
  AO22X1 U4608 ( .IN1(n4999), .IN2(n4294), .IN3(n5000), .IN4(n4295), .Q(n4971)
         );
  INVX0 U4609 ( .INP(n3064), .ZN(n4295) );
  AO222X1 U4610 ( .IN1(n4554), .IN2(n5355), .IN3(n4558), .IN4(n4556), .IN5(
        n4557), .IN6(n5367), .Q(n4524) );
  AO222X1 U4611 ( .IN1(n4583), .IN2(n5356), .IN3(n4587), .IN4(n4586), .IN5(
        n5368), .IN6(n4588), .Q(n4558) );
  AO222X1 U4612 ( .IN1(n4621), .IN2(n5357), .IN3(n4625), .IN4(n4591), .IN5(
        n4624), .IN6(n5369), .Q(n4587) );
  AO222X1 U4613 ( .IN1(n4654), .IN2(n5358), .IN3(n4656), .IN4(n4659), .IN5(
        n4658), .IN6(n5370), .Q(n4625) );
  AO222X1 U4614 ( .IN1(n4688), .IN2(n5359), .IN3(n4693), .IN4(n4691), .IN5(
        n4692), .IN6(n5371), .Q(n4659) );
  AO222X1 U4615 ( .IN1(n4724), .IN2(n5360), .IN3(n4728), .IN4(n4726), .IN5(
        n4727), .IN6(n5372), .Q(n4693) );
  AO222X1 U4616 ( .IN1(n4758), .IN2(n5361), .IN3(n4763), .IN4(n4761), .IN5(
        n4762), .IN6(n5373), .Q(n4728) );
  AO222X1 U4617 ( .IN1(n4797), .IN2(n5362), .IN3(n4800), .IN4(n4720), .IN5(
        n4753), .IN6(n5374), .Q(n4763) );
  AO222X1 U4618 ( .IN1(n4832), .IN2(n5363), .IN3(n4834), .IN4(n4837), .IN5(
        n4836), .IN6(n5375), .Q(n4800) );
  AO222X1 U4619 ( .IN1(n4876), .IN2(n5364), .IN3(n4881), .IN4(n4879), .IN5(
        n4880), .IN6(n5376), .Q(n4837) );
  AO222X1 U4620 ( .IN1(n4926), .IN2(n5365), .IN3(n4928), .IN4(n4931), .IN5(
        n4930), .IN6(n5377), .Q(n4881) );
  AO222X1 U4621 ( .IN1(n4970), .IN2(n5366), .IN3(n4975), .IN4(n4973), .IN5(
        n4974), .IN6(n5378), .Q(n4931) );
  AO22X1 U4622 ( .IN1(n4999), .IN2(n4293), .IN3(n5000), .IN4(n4294), .Q(n4975)
         );
  INVX0 U4623 ( .INP(n3065), .ZN(n4294) );
  AO222X1 U4624 ( .IN1(n5351), .IN2(n4522), .IN3(n4523), .IN4(n5099), .IN5(
        n4519), .IN6(n5101), .Q(n5093) );
  AO222X1 U4625 ( .IN1(n4554), .IN2(n5379), .IN3(n4557), .IN4(n5104), .IN5(
        n5367), .IN6(n4556), .Q(n5101) );
  NOR2X0 U4626 ( .IN1(n4523), .IN2(n4522), .QN(n4519) );
  AO222X1 U4627 ( .IN1(n4554), .IN2(n5104), .IN3(n4557), .IN4(n5102), .IN5(
        n5379), .IN6(n4556), .Q(n5099) );
  AO222X1 U4628 ( .IN1(n4583), .IN2(n5107), .IN3(n5105), .IN4(n4588), .IN5(
        n5380), .IN6(n4586), .Q(n5102) );
  AO222X1 U4629 ( .IN1(n4621), .IN2(n5110), .IN3(n4624), .IN4(n5108), .IN5(
        n5381), .IN6(n4591), .Q(n5105) );
  AO222X1 U4630 ( .IN1(n4654), .IN2(n5113), .IN3(n4658), .IN4(n5111), .IN5(
        n4656), .IN6(n5382), .Q(n5108) );
  AO222X1 U4631 ( .IN1(n4688), .IN2(n5116), .IN3(n4692), .IN4(n5114), .IN5(
        n5383), .IN6(n4691), .Q(n5111) );
  AO222X1 U4632 ( .IN1(n4724), .IN2(n5119), .IN3(n4727), .IN4(n5117), .IN5(
        n5384), .IN6(n4726), .Q(n5114) );
  AO222X1 U4633 ( .IN1(n4758), .IN2(n5122), .IN3(n4762), .IN4(n5120), .IN5(
        n5385), .IN6(n4761), .Q(n5117) );
  AO222X1 U4634 ( .IN1(n4797), .IN2(n5125), .IN3(n4753), .IN4(n5123), .IN5(
        n5386), .IN6(n4720), .Q(n5120) );
  AO222X1 U4635 ( .IN1(n4832), .IN2(n5128), .IN3(n4836), .IN4(n5126), .IN5(
        n4834), .IN6(n5387), .Q(n5123) );
  AO222X1 U4636 ( .IN1(n4876), .IN2(n5131), .IN3(n4880), .IN4(n5129), .IN5(
        n5388), .IN6(n4879), .Q(n5126) );
  AO222X1 U4637 ( .IN1(n4926), .IN2(n5134), .IN3(n4930), .IN4(n5132), .IN5(
        n4928), .IN6(n5389), .Q(n5129) );
  AO222X1 U4638 ( .IN1(n4970), .IN2(n5137), .IN3(n4974), .IN4(n5135), .IN5(
        n5390), .IN6(n4973), .Q(n5132) );
  AO22X1 U4639 ( .IN1(n4999), .IN2(n4266), .IN3(n5000), .IN4(n4267), .Q(n5135)
         );
  AO222X1 U4640 ( .IN1(n4583), .IN2(n5380), .IN3(n5107), .IN4(n4588), .IN5(
        n5391), .IN6(n4586), .Q(n5104) );
  AO222X1 U4641 ( .IN1(n4621), .IN2(n5381), .IN3(n4624), .IN4(n5110), .IN5(
        n5392), .IN6(n4591), .Q(n5107) );
  AO222X1 U4642 ( .IN1(n4654), .IN2(n5382), .IN3(n4658), .IN4(n5113), .IN5(
        n4656), .IN6(n5393), .Q(n5110) );
  AO222X1 U4643 ( .IN1(n4688), .IN2(n5383), .IN3(n4692), .IN4(n5116), .IN5(
        n5394), .IN6(n4691), .Q(n5113) );
  AO222X1 U4644 ( .IN1(n4724), .IN2(n5384), .IN3(n4727), .IN4(n5119), .IN5(
        n5395), .IN6(n4726), .Q(n5116) );
  AO222X1 U4645 ( .IN1(n4758), .IN2(n5385), .IN3(n4762), .IN4(n5122), .IN5(
        n5396), .IN6(n4761), .Q(n5119) );
  AO222X1 U4646 ( .IN1(n4797), .IN2(n5386), .IN3(n4753), .IN4(n5125), .IN5(
        n5397), .IN6(n4720), .Q(n5122) );
  AO222X1 U4647 ( .IN1(n4832), .IN2(n5387), .IN3(n4836), .IN4(n5128), .IN5(
        n4834), .IN6(n5398), .Q(n5125) );
  AO222X1 U4648 ( .IN1(n4876), .IN2(n5388), .IN3(n4880), .IN4(n5131), .IN5(
        n5399), .IN6(n4879), .Q(n5128) );
  AO222X1 U4649 ( .IN1(n4926), .IN2(n5389), .IN3(n4930), .IN4(n5134), .IN5(
        n4928), .IN6(n5400), .Q(n5131) );
  AO222X1 U4650 ( .IN1(n4970), .IN2(n5390), .IN3(n4974), .IN4(n5137), .IN5(
        n5401), .IN6(n4973), .Q(n5134) );
  AO22X1 U4651 ( .IN1(n4999), .IN2(n4267), .IN3(n5000), .IN4(n4268), .Q(n5137)
         );
  INVX0 U4652 ( .INP(n5017), .ZN(n4523) );
  AO21X1 U4653 ( .IN1(n5402), .IN2(n5403), .IN3(n5404), .Q(n5017) );
  NAND2X0 U4654 ( .IN1(n5405), .IN2(n5406), .QN(n5403) );
  AO21X1 U4655 ( .IN1(n5402), .IN2(n5407), .IN3(n5404), .Q(n4522) );
  AO21X1 U4656 ( .IN1(n5408), .IN2(n3803), .IN3(n5409), .Q(n5407) );
  AO222X1 U4657 ( .IN1(n4557), .IN2(n5379), .IN3(n5355), .IN4(n4556), .IN5(
        n4554), .IN6(n5367), .Q(n5351) );
  AO222X1 U4658 ( .IN1(n5391), .IN2(n4588), .IN3(n5368), .IN4(n4586), .IN5(
        n4583), .IN6(n5410), .Q(n5367) );
  NOR2X0 U4659 ( .IN1(n4556), .IN2(n4557), .QN(n4554) );
  NAND2X0 U4660 ( .IN1(n5310), .IN2(n5411), .QN(n4556) );
  NAND3X0 U4661 ( .IN1(\r150/A[3] ), .IN2(n5412), .IN3(n5402), .QN(n5411) );
  AO222X1 U4662 ( .IN1(n4583), .IN2(n5368), .IN3(n5356), .IN4(n4586), .IN5(
        n5410), .IN6(n4588), .Q(n5355) );
  AO222X1 U4663 ( .IN1(n4621), .IN2(n5369), .IN3(n5357), .IN4(n4591), .IN5(
        n4624), .IN6(n5413), .Q(n5356) );
  AO222X1 U4664 ( .IN1(n4654), .IN2(n5370), .IN3(n4656), .IN4(n5358), .IN5(
        n4658), .IN6(n5414), .Q(n5357) );
  AO222X1 U4665 ( .IN1(n4688), .IN2(n5371), .IN3(n5359), .IN4(n4691), .IN5(
        n4692), .IN6(n5415), .Q(n5358) );
  AO222X1 U4666 ( .IN1(n4724), .IN2(n5372), .IN3(n5360), .IN4(n4726), .IN5(
        n4727), .IN6(n5416), .Q(n5359) );
  AO222X1 U4667 ( .IN1(n4758), .IN2(n5373), .IN3(n5361), .IN4(n4761), .IN5(
        n4762), .IN6(n5417), .Q(n5360) );
  AO222X1 U4668 ( .IN1(n4797), .IN2(n5374), .IN3(n5362), .IN4(n4720), .IN5(
        n4753), .IN6(n5418), .Q(n5361) );
  AO222X1 U4669 ( .IN1(n4832), .IN2(n5375), .IN3(n4834), .IN4(n5363), .IN5(
        n4836), .IN6(n5419), .Q(n5362) );
  AO222X1 U4670 ( .IN1(n4876), .IN2(n5376), .IN3(n5364), .IN4(n4879), .IN5(
        n4880), .IN6(n5420), .Q(n5363) );
  AO222X1 U4671 ( .IN1(n4926), .IN2(n5377), .IN3(n4928), .IN4(n5365), .IN5(
        n4930), .IN6(n5421), .Q(n5364) );
  AO222X1 U4672 ( .IN1(n4970), .IN2(n5378), .IN3(n5366), .IN4(n4973), .IN5(
        n4974), .IN6(n5422), .Q(n5365) );
  AO22X1 U4673 ( .IN1(n4999), .IN2(n4292), .IN3(n5000), .IN4(n4293), .Q(n5366)
         );
  INVX0 U4674 ( .INP(n3066), .ZN(n4293) );
  AO222X1 U4675 ( .IN1(n4621), .IN2(n5413), .IN3(n5369), .IN4(n4591), .IN5(
        n4624), .IN6(n5423), .Q(n5368) );
  AO222X1 U4676 ( .IN1(n4654), .IN2(n5414), .IN3(n4656), .IN4(n5370), .IN5(
        n4658), .IN6(n5424), .Q(n5369) );
  AO222X1 U4677 ( .IN1(n4688), .IN2(n5415), .IN3(n5371), .IN4(n4691), .IN5(
        n4692), .IN6(n5425), .Q(n5370) );
  AO222X1 U4678 ( .IN1(n4724), .IN2(n5416), .IN3(n5372), .IN4(n4726), .IN5(
        n4727), .IN6(n5426), .Q(n5371) );
  AO222X1 U4679 ( .IN1(n4758), .IN2(n5417), .IN3(n5373), .IN4(n4761), .IN5(
        n4762), .IN6(n5427), .Q(n5372) );
  AO222X1 U4680 ( .IN1(n4797), .IN2(n5418), .IN3(n5374), .IN4(n4720), .IN5(
        n4753), .IN6(n5428), .Q(n5373) );
  AO222X1 U4681 ( .IN1(n4832), .IN2(n5419), .IN3(n4834), .IN4(n5375), .IN5(
        n4836), .IN6(n5429), .Q(n5374) );
  AO222X1 U4682 ( .IN1(n4876), .IN2(n5420), .IN3(n5376), .IN4(n4879), .IN5(
        n4880), .IN6(n5430), .Q(n5375) );
  AO222X1 U4683 ( .IN1(n4926), .IN2(n5421), .IN3(n4928), .IN4(n5377), .IN5(
        n4930), .IN6(n5431), .Q(n5376) );
  AO222X1 U4684 ( .IN1(n4970), .IN2(n5422), .IN3(n5378), .IN4(n4973), .IN5(
        n4974), .IN6(n5432), .Q(n5377) );
  AO22X1 U4685 ( .IN1(n4999), .IN2(n4291), .IN3(n5000), .IN4(n4292), .Q(n5378)
         );
  INVX0 U4686 ( .INP(n3067), .ZN(n4292) );
  AO222X1 U4687 ( .IN1(n5410), .IN2(n4586), .IN3(n5380), .IN4(n4588), .IN5(
        n4583), .IN6(n5391), .Q(n5379) );
  AO222X1 U4688 ( .IN1(n4621), .IN2(n5433), .IN3(n4624), .IN4(n5392), .IN5(
        n5423), .IN6(n4591), .Q(n5391) );
  NOR2X0 U4689 ( .IN1(n4586), .IN2(n4588), .QN(n4583) );
  INVX0 U4690 ( .INP(n4618), .ZN(n4588) );
  AO21X1 U4691 ( .IN1(n5434), .IN2(n5435), .IN3(n5436), .Q(n4618) );
  AO222X1 U4692 ( .IN1(n4621), .IN2(n5392), .IN3(n4624), .IN4(n5381), .IN5(
        n5433), .IN6(n4591), .Q(n5380) );
  AO222X1 U4693 ( .IN1(n4654), .IN2(n5393), .IN3(n4658), .IN4(n5382), .IN5(
        n4656), .IN6(n5437), .Q(n5381) );
  AO222X1 U4694 ( .IN1(n4688), .IN2(n5394), .IN3(n4692), .IN4(n5383), .IN5(
        n5438), .IN6(n4691), .Q(n5382) );
  AO222X1 U4695 ( .IN1(n4724), .IN2(n5395), .IN3(n4727), .IN4(n5384), .IN5(
        n5439), .IN6(n4726), .Q(n5383) );
  AO222X1 U4696 ( .IN1(n4758), .IN2(n5396), .IN3(n4762), .IN4(n5385), .IN5(
        n5440), .IN6(n4761), .Q(n5384) );
  AO222X1 U4697 ( .IN1(n4797), .IN2(n5397), .IN3(n4753), .IN4(n5386), .IN5(
        n5441), .IN6(n4720), .Q(n5385) );
  AO222X1 U4698 ( .IN1(n4832), .IN2(n5398), .IN3(n4836), .IN4(n5387), .IN5(
        n4834), .IN6(n5442), .Q(n5386) );
  AO222X1 U4699 ( .IN1(n4876), .IN2(n5399), .IN3(n4880), .IN4(n5388), .IN5(
        n5443), .IN6(n4879), .Q(n5387) );
  AO222X1 U4700 ( .IN1(n4926), .IN2(n5400), .IN3(n4930), .IN4(n5389), .IN5(
        n4928), .IN6(n5444), .Q(n5388) );
  AO222X1 U4701 ( .IN1(n4970), .IN2(n5401), .IN3(n4974), .IN4(n5390), .IN5(
        n5445), .IN6(n4973), .Q(n5389) );
  AO22X1 U4702 ( .IN1(n4999), .IN2(n4268), .IN3(n5000), .IN4(n4269), .Q(n5390)
         );
  AO222X1 U4703 ( .IN1(n4654), .IN2(n5437), .IN3(n4658), .IN4(n5393), .IN5(
        n4656), .IN6(n5446), .Q(n5392) );
  AO222X1 U4704 ( .IN1(n4688), .IN2(n5438), .IN3(n4692), .IN4(n5394), .IN5(
        n5447), .IN6(n4691), .Q(n5393) );
  AO222X1 U4705 ( .IN1(n4724), .IN2(n5439), .IN3(n4727), .IN4(n5395), .IN5(
        n5448), .IN6(n4726), .Q(n5394) );
  AO222X1 U4706 ( .IN1(n4758), .IN2(n5440), .IN3(n4762), .IN4(n5396), .IN5(
        n5449), .IN6(n4761), .Q(n5395) );
  AO222X1 U4707 ( .IN1(n4797), .IN2(n5441), .IN3(n4753), .IN4(n5397), .IN5(
        n5450), .IN6(n4720), .Q(n5396) );
  AO222X1 U4708 ( .IN1(n4832), .IN2(n5442), .IN3(n4836), .IN4(n5398), .IN5(
        n4834), .IN6(n5451), .Q(n5397) );
  AO222X1 U4709 ( .IN1(n4876), .IN2(n5443), .IN3(n4880), .IN4(n5399), .IN5(
        n5452), .IN6(n4879), .Q(n5398) );
  AO222X1 U4710 ( .IN1(n4926), .IN2(n5444), .IN3(n4930), .IN4(n5400), .IN5(
        n4928), .IN6(n5453), .Q(n5399) );
  AO222X1 U4711 ( .IN1(n4970), .IN2(n5445), .IN3(n4974), .IN4(n5401), .IN5(
        n5454), .IN6(n4973), .Q(n5400) );
  AO22X1 U4712 ( .IN1(n4999), .IN2(n4269), .IN3(n5000), .IN4(n4270), .Q(n5401)
         );
  INVX0 U4713 ( .INP(n5337), .ZN(n4586) );
  OA21X1 U4714 ( .IN1(n5455), .IN2(\r150/A[3] ), .IN3(n5456), .Q(n5337) );
  AO222X1 U4715 ( .IN1(n4624), .IN2(n5433), .IN3(n5413), .IN4(n4591), .IN5(
        n4621), .IN6(n5423), .Q(n5410) );
  AO222X1 U4716 ( .IN1(n4658), .IN2(n5446), .IN3(n4656), .IN4(n5424), .IN5(
        n4654), .IN6(n5457), .Q(n5423) );
  NOR2X0 U4717 ( .IN1(n4591), .IN2(n4624), .QN(n4621) );
  AO21X1 U4718 ( .IN1(n5458), .IN2(n5434), .IN3(n5459), .Q(n4591) );
  AO222X1 U4719 ( .IN1(n4654), .IN2(n5424), .IN3(n4656), .IN4(n5414), .IN5(
        n4658), .IN6(n5457), .Q(n5413) );
  AO222X1 U4720 ( .IN1(n4688), .IN2(n5425), .IN3(n5415), .IN4(n4691), .IN5(
        n4692), .IN6(n5460), .Q(n5414) );
  AO222X1 U4721 ( .IN1(n4724), .IN2(n5426), .IN3(n5416), .IN4(n4726), .IN5(
        n4727), .IN6(n5461), .Q(n5415) );
  AO222X1 U4722 ( .IN1(n4758), .IN2(n5427), .IN3(n5417), .IN4(n4761), .IN5(
        n4762), .IN6(n5462), .Q(n5416) );
  AO222X1 U4723 ( .IN1(n4797), .IN2(n5428), .IN3(n5418), .IN4(n4720), .IN5(
        n4753), .IN6(n5463), .Q(n5417) );
  AO222X1 U4724 ( .IN1(n4832), .IN2(n5429), .IN3(n4834), .IN4(n5419), .IN5(
        n4836), .IN6(n5464), .Q(n5418) );
  AO222X1 U4725 ( .IN1(n4876), .IN2(n5430), .IN3(n5420), .IN4(n4879), .IN5(
        n4880), .IN6(n5465), .Q(n5419) );
  AO222X1 U4726 ( .IN1(n4926), .IN2(n5431), .IN3(n4928), .IN4(n5421), .IN5(
        n4930), .IN6(n5466), .Q(n5420) );
  AO222X1 U4727 ( .IN1(n4970), .IN2(n5432), .IN3(n5422), .IN4(n4973), .IN5(
        n4974), .IN6(n5467), .Q(n5421) );
  AO22X1 U4728 ( .IN1(n4999), .IN2(n4290), .IN3(n5000), .IN4(n4291), .Q(n5422)
         );
  INVX0 U4729 ( .INP(n3068), .ZN(n4291) );
  AO222X1 U4730 ( .IN1(n4688), .IN2(n5460), .IN3(n5425), .IN4(n4691), .IN5(
        n4692), .IN6(n5468), .Q(n5424) );
  AO222X1 U4731 ( .IN1(n4724), .IN2(n5461), .IN3(n5426), .IN4(n4726), .IN5(
        n4727), .IN6(n5469), .Q(n5425) );
  AO222X1 U4732 ( .IN1(n4758), .IN2(n5462), .IN3(n5427), .IN4(n4761), .IN5(
        n4762), .IN6(n5470), .Q(n5426) );
  AO222X1 U4733 ( .IN1(n4797), .IN2(n5463), .IN3(n5428), .IN4(n4720), .IN5(
        n4753), .IN6(n5471), .Q(n5427) );
  AO222X1 U4734 ( .IN1(n4832), .IN2(n5464), .IN3(n4834), .IN4(n5429), .IN5(
        n4836), .IN6(n5472), .Q(n5428) );
  AO222X1 U4735 ( .IN1(n4876), .IN2(n5465), .IN3(n5430), .IN4(n4879), .IN5(
        n4880), .IN6(n5473), .Q(n5429) );
  AO222X1 U4736 ( .IN1(n4926), .IN2(n5466), .IN3(n4928), .IN4(n5431), .IN5(
        n4930), .IN6(n5474), .Q(n5430) );
  AO222X1 U4737 ( .IN1(n4970), .IN2(n5467), .IN3(n5432), .IN4(n4973), .IN5(
        n4974), .IN6(n5475), .Q(n5431) );
  AO22X1 U4738 ( .IN1(n4999), .IN2(n4289), .IN3(n5000), .IN4(n4290), .Q(n5432)
         );
  INVX0 U4739 ( .INP(n3069), .ZN(n4290) );
  AO222X1 U4740 ( .IN1(n4656), .IN2(n5457), .IN3(n4658), .IN4(n5437), .IN5(
        n4654), .IN6(n5446), .Q(n5433) );
  AO222X1 U4741 ( .IN1(n4688), .IN2(n5476), .IN3(n4692), .IN4(n5447), .IN5(
        n5468), .IN6(n4691), .Q(n5446) );
  NOR2X0 U4742 ( .IN1(n4651), .IN2(n4515), .QN(n4654) );
  AO222X1 U4743 ( .IN1(n4688), .IN2(n5447), .IN3(n4692), .IN4(n5438), .IN5(
        n5476), .IN6(n4691), .Q(n5437) );
  AO222X1 U4744 ( .IN1(n4724), .IN2(n5448), .IN3(n4727), .IN4(n5439), .IN5(
        n5477), .IN6(n4726), .Q(n5438) );
  AO222X1 U4745 ( .IN1(n4758), .IN2(n5449), .IN3(n4762), .IN4(n5440), .IN5(
        n5478), .IN6(n4761), .Q(n5439) );
  AO222X1 U4746 ( .IN1(n4797), .IN2(n5450), .IN3(n4753), .IN4(n5441), .IN5(
        n5479), .IN6(n4720), .Q(n5440) );
  AO222X1 U4747 ( .IN1(n4832), .IN2(n5451), .IN3(n4836), .IN4(n5442), .IN5(
        n4834), .IN6(n5480), .Q(n5441) );
  AO222X1 U4748 ( .IN1(n4876), .IN2(n5452), .IN3(n4880), .IN4(n5443), .IN5(
        n5481), .IN6(n4879), .Q(n5442) );
  AO222X1 U4749 ( .IN1(n4926), .IN2(n5453), .IN3(n4930), .IN4(n5444), .IN5(
        n4928), .IN6(n5482), .Q(n5443) );
  AO222X1 U4750 ( .IN1(n4970), .IN2(n5454), .IN3(n4974), .IN4(n5445), .IN5(
        n5483), .IN6(n4973), .Q(n5444) );
  AO22X1 U4751 ( .IN1(n4999), .IN2(n4270), .IN3(n5000), .IN4(n4271), .Q(n5445)
         );
  AO222X1 U4752 ( .IN1(n4724), .IN2(n5477), .IN3(n4727), .IN4(n5448), .IN5(
        n5484), .IN6(n4726), .Q(n5447) );
  AO222X1 U4753 ( .IN1(n4758), .IN2(n5478), .IN3(n4762), .IN4(n5449), .IN5(
        n5485), .IN6(n4761), .Q(n5448) );
  AO222X1 U4754 ( .IN1(n4797), .IN2(n5479), .IN3(n4753), .IN4(n5450), .IN5(
        n5486), .IN6(n4720), .Q(n5449) );
  AO222X1 U4755 ( .IN1(n4832), .IN2(n5480), .IN3(n4836), .IN4(n5451), .IN5(
        n4834), .IN6(n5487), .Q(n5450) );
  AO222X1 U4756 ( .IN1(n4876), .IN2(n5481), .IN3(n4880), .IN4(n5452), .IN5(
        n5488), .IN6(n4879), .Q(n5451) );
  AO222X1 U4757 ( .IN1(n4926), .IN2(n5482), .IN3(n4930), .IN4(n5453), .IN5(
        n4928), .IN6(n5489), .Q(n5452) );
  AO222X1 U4758 ( .IN1(n4970), .IN2(n5483), .IN3(n4974), .IN4(n5454), .IN5(
        n5490), .IN6(n4973), .Q(n5453) );
  AO22X1 U4759 ( .IN1(n4999), .IN2(n4271), .IN3(n5000), .IN4(n4272), .Q(n5454)
         );
  NOR2X0 U4760 ( .IN1(n5491), .IN2(n4651), .QN(n4658) );
  AO222X1 U4761 ( .IN1(n4692), .IN2(n5476), .IN3(n5460), .IN4(n4691), .IN5(
        n4688), .IN6(n5468), .Q(n5457) );
  AO222X1 U4762 ( .IN1(n4727), .IN2(n5484), .IN3(n5469), .IN4(n4726), .IN5(
        n4724), .IN6(n5492), .Q(n5468) );
  NOR2X0 U4763 ( .IN1(n4691), .IN2(n4692), .QN(n4688) );
  AO21X1 U4764 ( .IN1(n5458), .IN2(n5412), .IN3(n5436), .Q(n4691) );
  AOI21X1 U4765 ( .IN1(n5455), .IN2(n5310), .IN3(n5493), .QN(n5436) );
  AO222X1 U4766 ( .IN1(n4724), .IN2(n5469), .IN3(n5461), .IN4(n4726), .IN5(
        n4727), .IN6(n5492), .Q(n5460) );
  AO222X1 U4767 ( .IN1(n4758), .IN2(n5470), .IN3(n5462), .IN4(n4761), .IN5(
        n4762), .IN6(n5494), .Q(n5461) );
  AO222X1 U4768 ( .IN1(n4797), .IN2(n5471), .IN3(n5463), .IN4(n4720), .IN5(
        n4753), .IN6(n5495), .Q(n5462) );
  AO222X1 U4769 ( .IN1(n4832), .IN2(n5472), .IN3(n4834), .IN4(n5464), .IN5(
        n4836), .IN6(n5496), .Q(n5463) );
  AO222X1 U4770 ( .IN1(n4876), .IN2(n5473), .IN3(n5465), .IN4(n4879), .IN5(
        n4880), .IN6(n5497), .Q(n5464) );
  AO222X1 U4771 ( .IN1(n4926), .IN2(n5474), .IN3(n4928), .IN4(n5466), .IN5(
        n4930), .IN6(n5498), .Q(n5465) );
  AO222X1 U4772 ( .IN1(n4970), .IN2(n5475), .IN3(n5467), .IN4(n4973), .IN5(
        n4974), .IN6(n5499), .Q(n5466) );
  AO22X1 U4773 ( .IN1(n4999), .IN2(n4288), .IN3(n5000), .IN4(n4289), .Q(n5467)
         );
  INVX0 U4774 ( .INP(n3070), .ZN(n4289) );
  AO222X1 U4775 ( .IN1(n4758), .IN2(n5494), .IN3(n5470), .IN4(n4761), .IN5(
        n4762), .IN6(n5500), .Q(n5469) );
  AO222X1 U4776 ( .IN1(n4797), .IN2(n5495), .IN3(n5471), .IN4(n4720), .IN5(
        n4753), .IN6(n5501), .Q(n5470) );
  AO222X1 U4777 ( .IN1(n4832), .IN2(n5496), .IN3(n4834), .IN4(n5472), .IN5(
        n4836), .IN6(n5502), .Q(n5471) );
  AO222X1 U4778 ( .IN1(n4876), .IN2(n5497), .IN3(n5473), .IN4(n4879), .IN5(
        n4880), .IN6(n5503), .Q(n5472) );
  AO222X1 U4779 ( .IN1(n4926), .IN2(n5498), .IN3(n4928), .IN4(n5474), .IN5(
        n4930), .IN6(n5504), .Q(n5473) );
  AO222X1 U4780 ( .IN1(n4970), .IN2(n5499), .IN3(n5475), .IN4(n4973), .IN5(
        n4974), .IN6(n5505), .Q(n5474) );
  AO22X1 U4781 ( .IN1(n4999), .IN2(n4287), .IN3(n5000), .IN4(n4288), .Q(n5475)
         );
  INVX0 U4782 ( .INP(n3071), .ZN(n4288) );
  AO222X1 U4783 ( .IN1(n4724), .IN2(n5484), .IN3(n4727), .IN4(n5477), .IN5(
        n5492), .IN6(n4726), .Q(n5476) );
  AO222X1 U4784 ( .IN1(n4762), .IN2(n5506), .IN3(n5494), .IN4(n4761), .IN5(
        n4758), .IN6(n5500), .Q(n5492) );
  AO222X1 U4785 ( .IN1(n4797), .IN2(n5501), .IN3(n5495), .IN4(n4720), .IN5(
        n4753), .IN6(n5507), .Q(n5494) );
  AO222X1 U4786 ( .IN1(n4832), .IN2(n5502), .IN3(n4834), .IN4(n5496), .IN5(
        n4836), .IN6(n5508), .Q(n5495) );
  AO222X1 U4787 ( .IN1(n4876), .IN2(n5503), .IN3(n5497), .IN4(n4879), .IN5(
        n4880), .IN6(n5509), .Q(n5496) );
  AO222X1 U4788 ( .IN1(n4926), .IN2(n5504), .IN3(n4928), .IN4(n5498), .IN5(
        n4930), .IN6(n5510), .Q(n5497) );
  AO222X1 U4789 ( .IN1(n4970), .IN2(n5505), .IN3(n5499), .IN4(n4973), .IN5(
        n4974), .IN6(n5511), .Q(n5498) );
  AO22X1 U4790 ( .IN1(n4999), .IN2(n4286), .IN3(n5000), .IN4(n4287), .Q(n5499)
         );
  INVX0 U4791 ( .INP(n3072), .ZN(n4287) );
  AO222X1 U4792 ( .IN1(n4758), .IN2(n5485), .IN3(n4762), .IN4(n5478), .IN5(
        n5506), .IN6(n4761), .Q(n5477) );
  AO222X1 U4793 ( .IN1(n4797), .IN2(n5486), .IN3(n4753), .IN4(n5479), .IN5(
        n5512), .IN6(n4720), .Q(n5478) );
  AO222X1 U4794 ( .IN1(n4832), .IN2(n5487), .IN3(n4836), .IN4(n5480), .IN5(
        n4834), .IN6(n5513), .Q(n5479) );
  AO222X1 U4795 ( .IN1(n4876), .IN2(n5488), .IN3(n4880), .IN4(n5481), .IN5(
        n5514), .IN6(n4879), .Q(n5480) );
  AO222X1 U4796 ( .IN1(n4926), .IN2(n5489), .IN3(n4930), .IN4(n5482), .IN5(
        n4928), .IN6(n5515), .Q(n5481) );
  AO222X1 U4797 ( .IN1(n4970), .IN2(n5490), .IN3(n4974), .IN4(n5483), .IN5(
        n5516), .IN6(n4973), .Q(n5482) );
  AO22X1 U4798 ( .IN1(n4999), .IN2(n4272), .IN3(n5000), .IN4(n4273), .Q(n5483)
         );
  AO222X1 U4799 ( .IN1(n4758), .IN2(n5506), .IN3(n4762), .IN4(n5485), .IN5(
        n5500), .IN6(n4761), .Q(n5484) );
  AO222X1 U4800 ( .IN1(n4753), .IN2(n5517), .IN3(n5501), .IN4(n4720), .IN5(
        n4797), .IN6(n5507), .Q(n5500) );
  AO222X1 U4801 ( .IN1(n4832), .IN2(n5508), .IN3(n4834), .IN4(n5502), .IN5(
        n4836), .IN6(n5518), .Q(n5501) );
  AO222X1 U4802 ( .IN1(n4876), .IN2(n5509), .IN3(n5503), .IN4(n4879), .IN5(
        n4880), .IN6(n5519), .Q(n5502) );
  AO222X1 U4803 ( .IN1(n4926), .IN2(n5510), .IN3(n4928), .IN4(n5504), .IN5(
        n4930), .IN6(n5520), .Q(n5503) );
  AO222X1 U4804 ( .IN1(n4970), .IN2(n5511), .IN3(n5505), .IN4(n4973), .IN5(
        n4974), .IN6(n5521), .Q(n5504) );
  AO22X1 U4805 ( .IN1(n4999), .IN2(n4285), .IN3(n5000), .IN4(n4286), .Q(n5505)
         );
  INVX0 U4806 ( .INP(n3073), .ZN(n4286) );
  AO222X1 U4807 ( .IN1(n4797), .IN2(n5512), .IN3(n4753), .IN4(n5486), .IN5(
        n5517), .IN6(n4720), .Q(n5485) );
  AO222X1 U4808 ( .IN1(n4832), .IN2(n5513), .IN3(n4836), .IN4(n5487), .IN5(
        n4834), .IN6(n5522), .Q(n5486) );
  AO222X1 U4809 ( .IN1(n4876), .IN2(n5514), .IN3(n4880), .IN4(n5488), .IN5(
        n5523), .IN6(n4879), .Q(n5487) );
  AO222X1 U4810 ( .IN1(n4926), .IN2(n5515), .IN3(n4930), .IN4(n5489), .IN5(
        n4928), .IN6(n5524), .Q(n5488) );
  AO222X1 U4811 ( .IN1(n4970), .IN2(n5516), .IN3(n4974), .IN4(n5490), .IN5(
        n5525), .IN6(n4973), .Q(n5489) );
  AO22X1 U4812 ( .IN1(n4999), .IN2(n4273), .IN3(n5000), .IN4(n4274), .Q(n5490)
         );
  AO222X1 U4813 ( .IN1(n4797), .IN2(n5517), .IN3(n4753), .IN4(n5512), .IN5(
        n5507), .IN6(n4720), .Q(n5506) );
  AO222X1 U4814 ( .IN1(n4836), .IN2(n5526), .IN3(n4834), .IN4(n5508), .IN5(
        n4832), .IN6(n5518), .Q(n5507) );
  AO222X1 U4815 ( .IN1(n4876), .IN2(n5519), .IN3(n5509), .IN4(n4879), .IN5(
        n4880), .IN6(n5527), .Q(n5508) );
  AO222X1 U4816 ( .IN1(n4926), .IN2(n5520), .IN3(n4928), .IN4(n5510), .IN5(
        n4930), .IN6(n5528), .Q(n5509) );
  AO222X1 U4817 ( .IN1(n4970), .IN2(n5521), .IN3(n5511), .IN4(n4973), .IN5(
        n4974), .IN6(n5529), .Q(n5510) );
  AO22X1 U4818 ( .IN1(n4999), .IN2(n4284), .IN3(n5000), .IN4(n4285), .Q(n5511)
         );
  INVX0 U4819 ( .INP(n3074), .ZN(n4285) );
  AO222X1 U4820 ( .IN1(n4832), .IN2(n5522), .IN3(n4836), .IN4(n5513), .IN5(
        n4834), .IN6(n5526), .Q(n5512) );
  AO222X1 U4821 ( .IN1(n4876), .IN2(n5523), .IN3(n4880), .IN4(n5514), .IN5(
        n5530), .IN6(n4879), .Q(n5513) );
  AO222X1 U4822 ( .IN1(n4926), .IN2(n5524), .IN3(n4930), .IN4(n5515), .IN5(
        n4928), .IN6(n5531), .Q(n5514) );
  AO222X1 U4823 ( .IN1(n4970), .IN2(n5525), .IN3(n4974), .IN4(n5516), .IN5(
        n5532), .IN6(n4973), .Q(n5515) );
  AO22X1 U4824 ( .IN1(n4999), .IN2(n4274), .IN3(n5000), .IN4(n4275), .Q(n5516)
         );
  INVX0 U4825 ( .INP(n3085), .ZN(n4274) );
  AO222X1 U4826 ( .IN1(n4834), .IN2(n5518), .IN3(n4836), .IN4(n5522), .IN5(
        n4832), .IN6(n5526), .Q(n5517) );
  AO222X1 U4827 ( .IN1(n4876), .IN2(n5533), .IN3(n4880), .IN4(n5530), .IN5(
        n5527), .IN6(n4879), .Q(n5526) );
  XOR2X1 U4828 ( .IN1(n4649), .IN2(n4826), .Q(n4832) );
  AO222X1 U4829 ( .IN1(n4876), .IN2(n5530), .IN3(n4880), .IN4(n5523), .IN5(
        n5533), .IN6(n4879), .Q(n5522) );
  AO222X1 U4830 ( .IN1(n4926), .IN2(n5531), .IN3(n4930), .IN4(n5524), .IN5(
        n4928), .IN6(n5534), .Q(n5523) );
  AO222X1 U4831 ( .IN1(n4970), .IN2(n5532), .IN3(n4974), .IN4(n5525), .IN5(
        n5535), .IN6(n4973), .Q(n5524) );
  AO22X1 U4832 ( .IN1(n4999), .IN2(n4275), .IN3(n5000), .IN4(n4276), .Q(n5525)
         );
  INVX0 U4833 ( .INP(n3084), .ZN(n4275) );
  AO222X1 U4834 ( .IN1(n4926), .IN2(n5534), .IN3(n4930), .IN4(n5531), .IN5(
        n4928), .IN6(n5536), .Q(n5530) );
  AO222X1 U4835 ( .IN1(n4970), .IN2(n5535), .IN3(n4974), .IN4(n5532), .IN5(
        n5537), .IN6(n4973), .Q(n5531) );
  AO22X1 U4836 ( .IN1(n4999), .IN2(n4276), .IN3(n5000), .IN4(n4277), .Q(n5532)
         );
  INVX0 U4837 ( .INP(n3083), .ZN(n4276) );
  AND2X1 U4838 ( .IN1(n4826), .IN2(n4649), .Q(n4836) );
  AO222X1 U4839 ( .IN1(n4880), .IN2(n5533), .IN3(n5519), .IN4(n4879), .IN5(
        n4876), .IN6(n5527), .Q(n5518) );
  AO222X1 U4840 ( .IN1(n4930), .IN2(n5536), .IN3(n4928), .IN4(n5528), .IN5(
        n4926), .IN6(n5538), .Q(n5527) );
  NOR2X0 U4841 ( .IN1(n4879), .IN2(n4880), .QN(n4876) );
  NAND3X0 U4842 ( .IN1(n5539), .IN2(n5540), .IN3(n5493), .QN(n4879) );
  AO222X1 U4843 ( .IN1(n4926), .IN2(n5528), .IN3(n4928), .IN4(n5520), .IN5(
        n4930), .IN6(n5538), .Q(n5519) );
  AO222X1 U4844 ( .IN1(n4970), .IN2(n5529), .IN3(n5521), .IN4(n4973), .IN5(
        n4974), .IN6(n5541), .Q(n5520) );
  AO22X1 U4845 ( .IN1(n4999), .IN2(n4283), .IN3(n5000), .IN4(n4284), .Q(n5521)
         );
  INVX0 U4846 ( .INP(n3075), .ZN(n4284) );
  AO222X1 U4847 ( .IN1(n4970), .IN2(n5541), .IN3(n5529), .IN4(n4973), .IN5(
        n4974), .IN6(n5542), .Q(n5528) );
  AO22X1 U4848 ( .IN1(n4999), .IN2(n4282), .IN3(n5000), .IN4(n4283), .Q(n5529)
         );
  INVX0 U4849 ( .INP(n3076), .ZN(n4283) );
  AO222X1 U4850 ( .IN1(n4928), .IN2(n5538), .IN3(n4930), .IN4(n5534), .IN5(
        n4926), .IN6(n5536), .Q(n5533) );
  AO222X1 U4851 ( .IN1(n4970), .IN2(n5543), .IN3(n4974), .IN4(n5537), .IN5(
        n5542), .IN6(n4973), .Q(n5536) );
  XOR2X1 U4852 ( .IN1(n4916), .IN2(n4789), .Q(n4926) );
  AO222X1 U4853 ( .IN1(n4970), .IN2(n5537), .IN3(n4974), .IN4(n5535), .IN5(
        n5543), .IN6(n4973), .Q(n5534) );
  AO22X1 U4854 ( .IN1(n4999), .IN2(n4277), .IN3(n5000), .IN4(n4278), .Q(n5535)
         );
  INVX0 U4855 ( .INP(n3082), .ZN(n4277) );
  AO22X1 U4856 ( .IN1(n4999), .IN2(n4278), .IN3(n5000), .IN4(n4279), .Q(n5537)
         );
  INVX0 U4857 ( .INP(n3081), .ZN(n4278) );
  NOR2X0 U4858 ( .IN1(n5544), .IN2(n5545), .QN(n4930) );
  AO222X1 U4859 ( .IN1(n4974), .IN2(n5543), .IN3(n5541), .IN4(n4973), .IN5(
        n4970), .IN6(n5542), .Q(n5538) );
  AO22X1 U4860 ( .IN1(n4999), .IN2(n4280), .IN3(n5000), .IN4(n4281), .Q(n5542)
         );
  NOR2X0 U4861 ( .IN1(n4973), .IN2(n4974), .QN(n4970) );
  NAND4X0 U4862 ( .IN1(n5539), .IN2(n5546), .IN3(n5547), .IN4(n5548), .QN(
        n4973) );
  OA21X1 U4863 ( .IN1(n3803), .IN2(n5549), .IN3(n5550), .Q(n5548) );
  AO21X1 U4864 ( .IN1(n5551), .IN2(n5552), .IN3(n5553), .Q(n5547) );
  AO22X1 U4865 ( .IN1(n4999), .IN2(n4281), .IN3(n5000), .IN4(n4282), .Q(n5541)
         );
  INVX0 U4866 ( .INP(n3077), .ZN(n4282) );
  INVX0 U4867 ( .INP(n3078), .ZN(n4281) );
  AO22X1 U4868 ( .IN1(n4999), .IN2(n4279), .IN3(n5000), .IN4(n4280), .Q(n5543)
         );
  INVX0 U4869 ( .INP(n3079), .ZN(n4280) );
  NOR2X0 U4870 ( .IN1(n5001), .IN2(n4549), .QN(n5000) );
  INVX0 U4871 ( .INP(n3080), .ZN(n4279) );
  XOR2X1 U4872 ( .IN1(n4549), .IN2(n5001), .Q(n4999) );
  INVX0 U4873 ( .INP(n5341), .ZN(n5001) );
  NAND3X0 U4874 ( .IN1(n5554), .IN2(n5555), .IN3(n5493), .QN(n5341) );
  AND4X1 U4875 ( .IN1(n5556), .IN2(n5539), .IN3(n5310), .IN4(n5546), .Q(n4549)
         );
  AO21X1 U4876 ( .IN1(n3803), .IN2(n5353), .IN3(n5557), .Q(n5556) );
  INVX0 U4877 ( .INP(n5336), .ZN(n4974) );
  NAND3X0 U4878 ( .IN1(n5555), .IN2(n5406), .IN3(n5493), .QN(n5336) );
  NAND2X0 U4879 ( .IN1(\r150/A[3] ), .IN2(n5558), .QN(n5406) );
  NOR2X0 U4880 ( .IN1(n4916), .IN2(n4789), .QN(n4928) );
  INVX0 U4881 ( .INP(n5544), .ZN(n4789) );
  NAND4X0 U4882 ( .IN1(n5493), .IN2(n5559), .IN3(n5560), .IN4(n5539), .QN(
        n5544) );
  NAND2X0 U4883 ( .IN1(n5561), .IN2(n5558), .QN(n5560) );
  NAND2X0 U4884 ( .IN1(\r150/A[3] ), .IN2(n5562), .QN(n5559) );
  INVX0 U4885 ( .INP(n5545), .ZN(n4916) );
  NAND4X0 U4886 ( .IN1(n5493), .IN2(n5555), .IN3(n5563), .IN4(n5314), .QN(
        n5545) );
  OR2X1 U4887 ( .IN1(n5352), .IN2(n5551), .Q(n5563) );
  OA221X1 U4888 ( .IN1(n3803), .IN2(n5455), .IN3(n5549), .IN4(n5555), .IN5(
        n5493), .Q(n4880) );
  OA21X1 U4889 ( .IN1(n5314), .IN2(n5551), .IN3(n5555), .Q(n5455) );
  NOR2X0 U4890 ( .IN1(n4649), .IN2(n4826), .QN(n4834) );
  OA221X1 U4891 ( .IN1(n5313), .IN2(n5551), .IN3(n5555), .IN4(n5554), .IN5(
        n5493), .Q(n4826) );
  AND4X1 U4892 ( .IN1(n5550), .IN2(n5564), .IN3(n5565), .IN4(n5546), .Q(n4649)
         );
  NAND2X0 U4893 ( .IN1(n5566), .IN2(n5567), .QN(n5565) );
  NAND2X0 U4894 ( .IN1(n5568), .IN2(n5569), .QN(n5564) );
  NOR2X0 U4895 ( .IN1(n4720), .IN2(n4753), .QN(n4797) );
  NAND3X0 U4896 ( .IN1(n5570), .IN2(n5571), .IN3(n5572), .QN(n5163) );
  NAND2X0 U4897 ( .IN1(n5568), .IN2(n5566), .QN(n5570) );
  INVX0 U4898 ( .INP(n5539), .ZN(n5566) );
  INVX0 U4899 ( .INP(n5572), .ZN(n4720) );
  OA21X1 U4900 ( .IN1(n5539), .IN2(n5549), .IN3(n5493), .Q(n5572) );
  NAND2X0 U4901 ( .IN1(n5561), .IN2(\r150/A[3] ), .QN(n5539) );
  NOR2X0 U4902 ( .IN1(n4761), .IN2(n4762), .QN(n4758) );
  INVX0 U4903 ( .INP(n4919), .ZN(n4762) );
  NAND4X0 U4904 ( .IN1(n5493), .IN2(n5573), .IN3(n5571), .IN4(n5313), .QN(
        n4919) );
  NAND2X0 U4905 ( .IN1(n5561), .IN2(n5562), .QN(n5571) );
  NAND2X0 U4906 ( .IN1(n5434), .IN2(n3803), .QN(n5573) );
  OAI221X1 U4907 ( .IN1(n5313), .IN2(n5554), .IN3(n5314), .IN4(n5555), .IN5(
        n5493), .QN(n4761) );
  INVX0 U4908 ( .INP(n5561), .ZN(n5555) );
  NOR2X0 U4909 ( .IN1(n4726), .IN2(n4727), .QN(n4724) );
  AND4X1 U4910 ( .IN1(n5493), .IN2(n5574), .IN3(n5540), .IN4(n5313), .Q(n4727)
         );
  NAND3X0 U4911 ( .IN1(n5561), .IN2(n5575), .IN3(n5434), .QN(n5540) );
  NAND2X0 U4912 ( .IN1(n3803), .IN2(n5558), .QN(n5574) );
  NOR2X0 U4913 ( .IN1(n5569), .IN2(n5404), .QN(n5493) );
  NAND2X0 U4914 ( .IN1(n5354), .IN2(n5546), .QN(n4726) );
  OA21X1 U4915 ( .IN1(n5314), .IN2(n5353), .IN3(n5310), .Q(n5354) );
  INVX0 U4916 ( .INP(n5342), .ZN(n4692) );
  NAND3X0 U4917 ( .IN1(n5576), .IN2(n5313), .IN3(n5456), .QN(n5342) );
  AO21X1 U4918 ( .IN1(\r150/A[3] ), .IN2(n5553), .IN3(n5557), .Q(n5576) );
  INVX0 U4919 ( .INP(n5567), .ZN(n5557) );
  INVX0 U4920 ( .INP(n5569), .ZN(n5553) );
  NOR2X0 U4921 ( .IN1(n5550), .IN2(n4515), .QN(n4656) );
  INVX0 U4922 ( .INP(n5491), .ZN(n4515) );
  AO221X1 U4923 ( .IN1(n5402), .IN2(n5577), .IN3(n5458), .IN4(n5558), .IN5(
        n5404), .Q(n5491) );
  INVX0 U4924 ( .INP(n5578), .ZN(n5558) );
  INVX0 U4925 ( .INP(n5546), .ZN(n5458) );
  NAND2X0 U4926 ( .IN1(n5569), .IN2(\r150/A[3] ), .QN(n5546) );
  NAND2X0 U4927 ( .IN1(n5578), .IN2(n3803), .QN(n5577) );
  NOR2X0 U4928 ( .IN1(n5409), .IN2(n5568), .QN(n5578) );
  NOR2X0 U4929 ( .IN1(n5552), .IN2(n5551), .QN(n5568) );
  INVX0 U4930 ( .INP(n4651), .ZN(n5550) );
  AO21X1 U4931 ( .IN1(n5409), .IN2(n5569), .IN3(n5459), .Q(n4651) );
  INVX0 U4932 ( .INP(n4965), .ZN(n4624) );
  NAND4X0 U4933 ( .IN1(n5456), .IN2(n5579), .IN3(n5313), .IN4(n5352), .QN(
        n4965) );
  NAND2X0 U4934 ( .IN1(n5409), .IN2(n3803), .QN(n5352) );
  NAND2X0 U4935 ( .IN1(n5561), .IN2(n3803), .QN(n5313) );
  NAND2X0 U4936 ( .IN1(n5569), .IN2(n5562), .QN(n5579) );
  NOR2X0 U4937 ( .IN1(n5459), .IN2(n5435), .QN(n5456) );
  NAND2X0 U4938 ( .IN1(n5353), .IN2(n5310), .QN(n5459) );
  AOI221X1 U4939 ( .IN1(n5435), .IN2(n5562), .IN3(n5402), .IN4(n5567), .IN5(
        n5580), .QN(n4557) );
  NAND2X0 U4940 ( .IN1(n5554), .IN2(n5551), .QN(n5567) );
  INVX0 U4941 ( .INP(n5412), .ZN(n5554) );
  INVX0 U4942 ( .INP(n4685), .ZN(n4489) );
  AO221X1 U4943 ( .IN1(n5435), .IN2(n5412), .IN3(n5402), .IN4(n5562), .IN5(
        n5580), .Q(n4685) );
  AO21X1 U4944 ( .IN1(n5402), .IN2(n3803), .IN3(n5404), .Q(n5580) );
  INVX0 U4945 ( .INP(n5310), .ZN(n5404) );
  NAND2X0 U4946 ( .IN1(n3803), .IN2(n5344), .QN(n5310) );
  NAND3X0 U4947 ( .IN1(n3088), .IN2(n3087), .IN3(n3089), .QN(n5344) );
  INVX0 U4948 ( .INP(n5405), .ZN(n5562) );
  OA21X1 U4949 ( .IN1(n5549), .IN2(n5551), .IN3(n5314), .Q(n5405) );
  INVX0 U4950 ( .INP(n5575), .ZN(n5551) );
  NAND2X0 U4951 ( .IN1(n5549), .IN2(n5552), .QN(n5412) );
  INVX0 U4952 ( .INP(n5408), .ZN(n5552) );
  INVX0 U4953 ( .INP(n5409), .ZN(n5549) );
  INVX0 U4954 ( .INP(n5311), .ZN(n5435) );
  NAND2X0 U4955 ( .IN1(n5569), .IN2(n3803), .QN(n5311) );
  AND2X1 U4956 ( .IN1(n5089), .IN2(n5345), .Q(n4459) );
  AND3X1 U4957 ( .IN1(n5723), .IN2(n4415), .IN3(n5350), .Q(n5345) );
  INVX0 U4958 ( .INP(n4417), .ZN(n4415) );
  NOR3X0 U4959 ( .IN1(n4375), .IN2(n4408), .IN3(n4371), .QN(n4417) );
  NAND3X0 U4960 ( .IN1(n2991), .IN2(n2988), .IN3(n2994), .QN(n4408) );
  INVX0 U4961 ( .INP(n5343), .ZN(n5089) );
  NAND3X0 U4962 ( .IN1(n5575), .IN2(n5402), .IN3(n5434), .QN(n5343) );
  INVX0 U4963 ( .INP(n5314), .ZN(n5434) );
  NAND2X0 U4964 ( .IN1(n5408), .IN2(n5409), .QN(n5314) );
  MUX21X1 U4965 ( .IN1(n4267), .IN2(n4381), .S(\r150/A[3] ), .Q(n5409) );
  MUX21X1 U4966 ( .IN1(n4266), .IN2(n4383), .S(\r150/A[3] ), .Q(n5408) );
  INVX0 U4967 ( .INP(n5353), .ZN(n5402) );
  NAND2X0 U4968 ( .IN1(n5561), .IN2(n5569), .QN(n5353) );
  MUX21X1 U4969 ( .IN1(n4269), .IN2(n4371), .S(\r150/A[3] ), .Q(n5569) );
  MUX21X1 U4970 ( .IN1(n4268), .IN2(n4375), .S(\r150/A[3] ), .Q(n5561) );
  MUX21X1 U4971 ( .IN1(n4265), .IN2(n4384), .S(\r150/A[3] ), .Q(n5575) );
  AND4X1 U4972 ( .IN1(n5581), .IN2(n5723), .IN3(n3844), .IN4(n3803), .Q(n4466)
         );
  AO221X1 U4973 ( .IN1(N3756), .IN2(n4473), .IN3(N3588), .IN4(n4465), .IN5(
        n5582), .Q(n5061) );
  AO222X1 U4974 ( .IN1(N3654), .IN2(n4505), .IN3(N3687), .IN4(n4471), .IN5(
        N3790), .IN6(n4474), .Q(n5582) );
  INVX0 U4975 ( .INP(n5044), .ZN(n4474) );
  NAND2X0 U4976 ( .IN1(n4410), .IN2(n3844), .QN(n5044) );
  INVX0 U4977 ( .INP(n5042), .ZN(n4410) );
  AND2X1 U4978 ( .IN1(n5583), .IN2(n3804), .Q(n4471) );
  AO22X1 U4979 ( .IN1(n4425), .IN2(n4406), .IN3(n5720), .IN4(n4407), .Q(n5583)
         );
  NOR2X0 U4980 ( .IN1(n3805), .IN2(n3843), .QN(n4407) );
  NOR3X0 U4981 ( .IN1(n4429), .IN2(n5724), .IN3(n5074), .QN(n4505) );
  AOI21X1 U4982 ( .IN1(n3804), .IN2(n5584), .IN3(n5074), .QN(n4465) );
  NAND2X0 U4983 ( .IN1(n4406), .IN2(n5724), .QN(n5584) );
  AND4X1 U4984 ( .IN1(n5581), .IN2(n4425), .IN3(n5585), .IN4(n3805), .Q(n4473)
         );
  NOR2X0 U4985 ( .IN1(n5720), .IN2(n5722), .QN(n5585) );
  INVX0 U4986 ( .INP(n5056), .ZN(n4425) );
  AND3X1 U4987 ( .IN1(n3088), .IN2(n3087), .IN3(n5586), .Q(n5581) );
  OA22X1 U4988 ( .IN1(n3089), .IN2(n3090), .IN3(n5587), .IN4(n3089), .Q(n5586)
         );
  NOR4X0 U4989 ( .IN1(n4268), .IN2(n4267), .IN3(n4266), .IN4(n4265), .QN(n5587) );
  MUX21X1 U4990 ( .IN1(\R[7][31] ), .IN2(n5588), .S(n5589), .Q(n3427) );
  MUX21X1 U4991 ( .IN1(\R[7][30] ), .IN2(n5590), .S(n5589), .Q(n3426) );
  MUX21X1 U4992 ( .IN1(\R[7][29] ), .IN2(n5591), .S(n5589), .Q(n3425) );
  MUX21X1 U4993 ( .IN1(\R[7][28] ), .IN2(n5592), .S(n5589), .Q(n3424) );
  MUX21X1 U4994 ( .IN1(\R[7][27] ), .IN2(n5593), .S(n5589), .Q(n3423) );
  MUX21X1 U4995 ( .IN1(\R[7][26] ), .IN2(n5594), .S(n5589), .Q(n3422) );
  MUX21X1 U4996 ( .IN1(\R[7][25] ), .IN2(n5595), .S(n5589), .Q(n3421) );
  MUX21X1 U4997 ( .IN1(\R[7][24] ), .IN2(n5596), .S(n5589), .Q(n3420) );
  MUX21X1 U4998 ( .IN1(\R[7][23] ), .IN2(n5597), .S(n5589), .Q(n3419) );
  MUX21X1 U4999 ( .IN1(\R[7][22] ), .IN2(n5598), .S(n5589), .Q(n3418) );
  MUX21X1 U5000 ( .IN1(\R[7][21] ), .IN2(n5599), .S(n5589), .Q(n3417) );
  MUX21X1 U5001 ( .IN1(\R[7][20] ), .IN2(n5600), .S(n5589), .Q(n3416) );
  MUX21X1 U5002 ( .IN1(\R[7][19] ), .IN2(n5601), .S(n5589), .Q(n3415) );
  MUX21X1 U5003 ( .IN1(\R[7][18] ), .IN2(n5602), .S(n5589), .Q(n3414) );
  MUX21X1 U5004 ( .IN1(\R[7][17] ), .IN2(n5603), .S(n5589), .Q(n3413) );
  MUX21X1 U5005 ( .IN1(\R[7][16] ), .IN2(n5604), .S(n5589), .Q(n3412) );
  MUX21X1 U5006 ( .IN1(\R[7][15] ), .IN2(n5605), .S(n5589), .Q(n3411) );
  MUX21X1 U5007 ( .IN1(\R[7][14] ), .IN2(n5606), .S(n5589), .Q(n3410) );
  MUX21X1 U5008 ( .IN1(\R[7][13] ), .IN2(n5607), .S(n5589), .Q(n3409) );
  MUX21X1 U5009 ( .IN1(\R[7][12] ), .IN2(n5608), .S(n5589), .Q(n3408) );
  MUX21X1 U5010 ( .IN1(\R[7][11] ), .IN2(n5609), .S(n5589), .Q(n3407) );
  MUX21X1 U5011 ( .IN1(\R[7][10] ), .IN2(n5610), .S(n5589), .Q(n3406) );
  MUX21X1 U5012 ( .IN1(\R[7][9] ), .IN2(n5611), .S(n5589), .Q(n3405) );
  MUX21X1 U5013 ( .IN1(\R[7][8] ), .IN2(n5612), .S(n5589), .Q(n3404) );
  MUX21X1 U5014 ( .IN1(\R[7][7] ), .IN2(n5613), .S(n5589), .Q(n3403) );
  MUX21X1 U5015 ( .IN1(\R[7][6] ), .IN2(n5614), .S(n5589), .Q(n3402) );
  MUX21X1 U5016 ( .IN1(\R[7][5] ), .IN2(n5615), .S(n5589), .Q(n3401) );
  MUX21X1 U5017 ( .IN1(\R[7][4] ), .IN2(n5616), .S(n5589), .Q(n3400) );
  MUX21X1 U5018 ( .IN1(\R[7][3] ), .IN2(n5617), .S(n5589), .Q(n3399) );
  MUX21X1 U5019 ( .IN1(\R[7][2] ), .IN2(n5618), .S(n5589), .Q(n3398) );
  MUX21X1 U5020 ( .IN1(\R[7][1] ), .IN2(n5619), .S(n5589), .Q(n3397) );
  MUX21X1 U5021 ( .IN1(\R[7][0] ), .IN2(n5620), .S(n5589), .Q(n3396) );
  AND3X1 U5022 ( .IN1(n3808), .IN2(n3806), .IN3(n5621), .Q(n5589) );
  MUX21X1 U5023 ( .IN1(\R[6][31] ), .IN2(n5588), .S(n5622), .Q(n3395) );
  MUX21X1 U5024 ( .IN1(\R[6][30] ), .IN2(n5590), .S(n5622), .Q(n3394) );
  MUX21X1 U5025 ( .IN1(\R[6][29] ), .IN2(n5591), .S(n5622), .Q(n3393) );
  MUX21X1 U5026 ( .IN1(\R[6][28] ), .IN2(n5592), .S(n5622), .Q(n3392) );
  MUX21X1 U5027 ( .IN1(\R[6][27] ), .IN2(n5593), .S(n5622), .Q(n3391) );
  MUX21X1 U5028 ( .IN1(\R[6][26] ), .IN2(n5594), .S(n5622), .Q(n3390) );
  MUX21X1 U5029 ( .IN1(\R[6][25] ), .IN2(n5595), .S(n5622), .Q(n3389) );
  MUX21X1 U5030 ( .IN1(\R[6][24] ), .IN2(n5596), .S(n5622), .Q(n3388) );
  MUX21X1 U5031 ( .IN1(\R[6][23] ), .IN2(n5597), .S(n5622), .Q(n3387) );
  MUX21X1 U5032 ( .IN1(\R[6][22] ), .IN2(n5598), .S(n5622), .Q(n3386) );
  MUX21X1 U5033 ( .IN1(\R[6][21] ), .IN2(n5599), .S(n5622), .Q(n3385) );
  MUX21X1 U5034 ( .IN1(\R[6][20] ), .IN2(n5600), .S(n5622), .Q(n3384) );
  MUX21X1 U5035 ( .IN1(\R[6][19] ), .IN2(n5601), .S(n5622), .Q(n3383) );
  MUX21X1 U5036 ( .IN1(\R[6][18] ), .IN2(n5602), .S(n5622), .Q(n3382) );
  MUX21X1 U5037 ( .IN1(\R[6][17] ), .IN2(n5603), .S(n5622), .Q(n3381) );
  MUX21X1 U5038 ( .IN1(\R[6][16] ), .IN2(n5604), .S(n5622), .Q(n3380) );
  MUX21X1 U5039 ( .IN1(\R[6][15] ), .IN2(n5605), .S(n5622), .Q(n3379) );
  MUX21X1 U5040 ( .IN1(\R[6][14] ), .IN2(n5606), .S(n5622), .Q(n3378) );
  MUX21X1 U5041 ( .IN1(\R[6][13] ), .IN2(n5607), .S(n5622), .Q(n3377) );
  MUX21X1 U5042 ( .IN1(\R[6][12] ), .IN2(n5608), .S(n5622), .Q(n3376) );
  MUX21X1 U5043 ( .IN1(\R[6][11] ), .IN2(n5609), .S(n5622), .Q(n3375) );
  MUX21X1 U5044 ( .IN1(\R[6][10] ), .IN2(n5610), .S(n5622), .Q(n3374) );
  MUX21X1 U5045 ( .IN1(\R[6][9] ), .IN2(n5611), .S(n5622), .Q(n3373) );
  MUX21X1 U5046 ( .IN1(\R[6][8] ), .IN2(n5612), .S(n5622), .Q(n3372) );
  MUX21X1 U5047 ( .IN1(\R[6][7] ), .IN2(n5613), .S(n5622), .Q(n3371) );
  MUX21X1 U5048 ( .IN1(\R[6][6] ), .IN2(n5614), .S(n5622), .Q(n3370) );
  MUX21X1 U5049 ( .IN1(\R[6][5] ), .IN2(n5615), .S(n5622), .Q(n3369) );
  MUX21X1 U5050 ( .IN1(\R[6][4] ), .IN2(n5616), .S(n5622), .Q(n3368) );
  MUX21X1 U5051 ( .IN1(\R[6][3] ), .IN2(n5617), .S(n5622), .Q(n3367) );
  MUX21X1 U5052 ( .IN1(\R[6][2] ), .IN2(n5618), .S(n5622), .Q(n3366) );
  MUX21X1 U5053 ( .IN1(\R[6][1] ), .IN2(n5619), .S(n5622), .Q(n3365) );
  MUX21X1 U5054 ( .IN1(\R[6][0] ), .IN2(n5620), .S(n5622), .Q(n3364) );
  AND3X1 U5055 ( .IN1(n3808), .IN2(n3806), .IN3(n5623), .Q(n5622) );
  MUX21X1 U5056 ( .IN1(\R[5][31] ), .IN2(n5588), .S(n5624), .Q(n3363) );
  MUX21X1 U5057 ( .IN1(\R[5][30] ), .IN2(n5590), .S(n5624), .Q(n3362) );
  MUX21X1 U5058 ( .IN1(\R[5][29] ), .IN2(n5591), .S(n5624), .Q(n3361) );
  MUX21X1 U5059 ( .IN1(\R[5][28] ), .IN2(n5592), .S(n5624), .Q(n3360) );
  MUX21X1 U5060 ( .IN1(\R[5][27] ), .IN2(n5593), .S(n5624), .Q(n3359) );
  MUX21X1 U5061 ( .IN1(\R[5][26] ), .IN2(n5594), .S(n5624), .Q(n3358) );
  MUX21X1 U5062 ( .IN1(\R[5][25] ), .IN2(n5595), .S(n5624), .Q(n3357) );
  MUX21X1 U5063 ( .IN1(\R[5][24] ), .IN2(n5596), .S(n5624), .Q(n3356) );
  MUX21X1 U5064 ( .IN1(\R[5][23] ), .IN2(n5597), .S(n5624), .Q(n3355) );
  MUX21X1 U5065 ( .IN1(\R[5][22] ), .IN2(n5598), .S(n5624), .Q(n3354) );
  MUX21X1 U5066 ( .IN1(\R[5][21] ), .IN2(n5599), .S(n5624), .Q(n3353) );
  MUX21X1 U5067 ( .IN1(\R[5][20] ), .IN2(n5600), .S(n5624), .Q(n3352) );
  MUX21X1 U5068 ( .IN1(\R[5][19] ), .IN2(n5601), .S(n5624), .Q(n3351) );
  MUX21X1 U5069 ( .IN1(\R[5][18] ), .IN2(n5602), .S(n5624), .Q(n3350) );
  MUX21X1 U5070 ( .IN1(\R[5][17] ), .IN2(n5603), .S(n5624), .Q(n3349) );
  MUX21X1 U5071 ( .IN1(\R[5][16] ), .IN2(n5604), .S(n5624), .Q(n3348) );
  MUX21X1 U5072 ( .IN1(\R[5][15] ), .IN2(n5605), .S(n5624), .Q(n3347) );
  MUX21X1 U5073 ( .IN1(\R[5][14] ), .IN2(n5606), .S(n5624), .Q(n3346) );
  MUX21X1 U5074 ( .IN1(\R[5][13] ), .IN2(n5607), .S(n5624), .Q(n3345) );
  MUX21X1 U5075 ( .IN1(\R[5][12] ), .IN2(n5608), .S(n5624), .Q(n3344) );
  MUX21X1 U5076 ( .IN1(\R[5][11] ), .IN2(n5609), .S(n5624), .Q(n3343) );
  MUX21X1 U5077 ( .IN1(\R[5][10] ), .IN2(n5610), .S(n5624), .Q(n3342) );
  MUX21X1 U5078 ( .IN1(\R[5][9] ), .IN2(n5611), .S(n5624), .Q(n3341) );
  MUX21X1 U5079 ( .IN1(\R[5][8] ), .IN2(n5612), .S(n5624), .Q(n3340) );
  MUX21X1 U5080 ( .IN1(\R[5][7] ), .IN2(n5613), .S(n5624), .Q(n3339) );
  MUX21X1 U5081 ( .IN1(\R[5][6] ), .IN2(n5614), .S(n5624), .Q(n3338) );
  MUX21X1 U5082 ( .IN1(\R[5][5] ), .IN2(n5615), .S(n5624), .Q(n3337) );
  MUX21X1 U5083 ( .IN1(\R[5][4] ), .IN2(n5616), .S(n5624), .Q(n3336) );
  MUX21X1 U5084 ( .IN1(\R[5][3] ), .IN2(n5617), .S(n5624), .Q(n3335) );
  MUX21X1 U5085 ( .IN1(\R[5][2] ), .IN2(n5618), .S(n5624), .Q(n3334) );
  MUX21X1 U5086 ( .IN1(\R[5][1] ), .IN2(n5619), .S(n5624), .Q(n3333) );
  MUX21X1 U5087 ( .IN1(\R[5][0] ), .IN2(n5620), .S(n5624), .Q(n3332) );
  AND3X1 U5088 ( .IN1(n5621), .IN2(n3808), .IN3(n5716), .Q(n5624) );
  MUX21X1 U5089 ( .IN1(\R[4][31] ), .IN2(n5588), .S(n5625), .Q(n3331) );
  MUX21X1 U5090 ( .IN1(\R[4][30] ), .IN2(n5590), .S(n5625), .Q(n3330) );
  MUX21X1 U5091 ( .IN1(\R[4][29] ), .IN2(n5591), .S(n5625), .Q(n3329) );
  MUX21X1 U5092 ( .IN1(\R[4][28] ), .IN2(n5592), .S(n5625), .Q(n3328) );
  MUX21X1 U5093 ( .IN1(\R[4][27] ), .IN2(n5593), .S(n5625), .Q(n3327) );
  MUX21X1 U5094 ( .IN1(\R[4][26] ), .IN2(n5594), .S(n5625), .Q(n3326) );
  MUX21X1 U5095 ( .IN1(\R[4][25] ), .IN2(n5595), .S(n5625), .Q(n3325) );
  MUX21X1 U5096 ( .IN1(\R[4][24] ), .IN2(n5596), .S(n5625), .Q(n3324) );
  MUX21X1 U5097 ( .IN1(\R[4][23] ), .IN2(n5597), .S(n5625), .Q(n3323) );
  MUX21X1 U5098 ( .IN1(\R[4][22] ), .IN2(n5598), .S(n5625), .Q(n3322) );
  MUX21X1 U5099 ( .IN1(\R[4][21] ), .IN2(n5599), .S(n5625), .Q(n3321) );
  MUX21X1 U5100 ( .IN1(\R[4][20] ), .IN2(n5600), .S(n5625), .Q(n3320) );
  MUX21X1 U5101 ( .IN1(\R[4][19] ), .IN2(n5601), .S(n5625), .Q(n3319) );
  MUX21X1 U5102 ( .IN1(\R[4][18] ), .IN2(n5602), .S(n5625), .Q(n3318) );
  MUX21X1 U5103 ( .IN1(\R[4][17] ), .IN2(n5603), .S(n5625), .Q(n3317) );
  MUX21X1 U5104 ( .IN1(\R[4][16] ), .IN2(n5604), .S(n5625), .Q(n3316) );
  MUX21X1 U5105 ( .IN1(\R[4][15] ), .IN2(n5605), .S(n5625), .Q(n3315) );
  MUX21X1 U5106 ( .IN1(\R[4][14] ), .IN2(n5606), .S(n5625), .Q(n3314) );
  MUX21X1 U5107 ( .IN1(\R[4][13] ), .IN2(n5607), .S(n5625), .Q(n3313) );
  MUX21X1 U5108 ( .IN1(\R[4][12] ), .IN2(n5608), .S(n5625), .Q(n3312) );
  MUX21X1 U5109 ( .IN1(\R[4][11] ), .IN2(n5609), .S(n5625), .Q(n3311) );
  MUX21X1 U5110 ( .IN1(\R[4][10] ), .IN2(n5610), .S(n5625), .Q(n3310) );
  MUX21X1 U5111 ( .IN1(\R[4][9] ), .IN2(n5611), .S(n5625), .Q(n3309) );
  MUX21X1 U5112 ( .IN1(\R[4][8] ), .IN2(n5612), .S(n5625), .Q(n3308) );
  MUX21X1 U5113 ( .IN1(\R[4][7] ), .IN2(n5613), .S(n5625), .Q(n3307) );
  MUX21X1 U5114 ( .IN1(\R[4][6] ), .IN2(n5614), .S(n5625), .Q(n3306) );
  MUX21X1 U5115 ( .IN1(\R[4][5] ), .IN2(n5615), .S(n5625), .Q(n3305) );
  MUX21X1 U5116 ( .IN1(\R[4][4] ), .IN2(n5616), .S(n5625), .Q(n3304) );
  MUX21X1 U5117 ( .IN1(\R[4][3] ), .IN2(n5617), .S(n5625), .Q(n3303) );
  MUX21X1 U5118 ( .IN1(\R[4][2] ), .IN2(n5618), .S(n5625), .Q(n3302) );
  MUX21X1 U5119 ( .IN1(\R[4][1] ), .IN2(n5619), .S(n5625), .Q(n3301) );
  MUX21X1 U5120 ( .IN1(\R[4][0] ), .IN2(n5620), .S(n5625), .Q(n3300) );
  AND3X1 U5121 ( .IN1(n5623), .IN2(n3808), .IN3(n5716), .Q(n5625) );
  MUX21X1 U5122 ( .IN1(\R[3][31] ), .IN2(n5588), .S(n5626), .Q(n3299) );
  MUX21X1 U5123 ( .IN1(\R[3][30] ), .IN2(n5590), .S(n5626), .Q(n3298) );
  MUX21X1 U5124 ( .IN1(\R[3][29] ), .IN2(n5591), .S(n5626), .Q(n3297) );
  MUX21X1 U5125 ( .IN1(\R[3][28] ), .IN2(n5592), .S(n5626), .Q(n3296) );
  MUX21X1 U5126 ( .IN1(\R[3][27] ), .IN2(n5593), .S(n5626), .Q(n3295) );
  MUX21X1 U5127 ( .IN1(\R[3][26] ), .IN2(n5594), .S(n5626), .Q(n3294) );
  MUX21X1 U5128 ( .IN1(\R[3][25] ), .IN2(n5595), .S(n5626), .Q(n3293) );
  MUX21X1 U5129 ( .IN1(\R[3][24] ), .IN2(n5596), .S(n5626), .Q(n3292) );
  MUX21X1 U5130 ( .IN1(\R[3][23] ), .IN2(n5597), .S(n5626), .Q(n3291) );
  MUX21X1 U5131 ( .IN1(\R[3][22] ), .IN2(n5598), .S(n5626), .Q(n3290) );
  MUX21X1 U5132 ( .IN1(\R[3][21] ), .IN2(n5599), .S(n5626), .Q(n3289) );
  MUX21X1 U5133 ( .IN1(\R[3][20] ), .IN2(n5600), .S(n5626), .Q(n3288) );
  MUX21X1 U5134 ( .IN1(\R[3][19] ), .IN2(n5601), .S(n5626), .Q(n3287) );
  MUX21X1 U5135 ( .IN1(\R[3][18] ), .IN2(n5602), .S(n5626), .Q(n3286) );
  MUX21X1 U5136 ( .IN1(\R[3][17] ), .IN2(n5603), .S(n5626), .Q(n3285) );
  MUX21X1 U5137 ( .IN1(\R[3][16] ), .IN2(n5604), .S(n5626), .Q(n3284) );
  MUX21X1 U5138 ( .IN1(\R[3][15] ), .IN2(n5605), .S(n5626), .Q(n3283) );
  MUX21X1 U5139 ( .IN1(\R[3][14] ), .IN2(n5606), .S(n5626), .Q(n3282) );
  MUX21X1 U5140 ( .IN1(\R[3][13] ), .IN2(n5607), .S(n5626), .Q(n3281) );
  MUX21X1 U5141 ( .IN1(\R[3][12] ), .IN2(n5608), .S(n5626), .Q(n3280) );
  MUX21X1 U5142 ( .IN1(\R[3][11] ), .IN2(n5609), .S(n5626), .Q(n3279) );
  MUX21X1 U5143 ( .IN1(\R[3][10] ), .IN2(n5610), .S(n5626), .Q(n3278) );
  MUX21X1 U5144 ( .IN1(\R[3][9] ), .IN2(n5611), .S(n5626), .Q(n3277) );
  MUX21X1 U5145 ( .IN1(\R[3][8] ), .IN2(n5612), .S(n5626), .Q(n3276) );
  MUX21X1 U5146 ( .IN1(\R[3][7] ), .IN2(n5613), .S(n5626), .Q(n3275) );
  MUX21X1 U5147 ( .IN1(\R[3][6] ), .IN2(n5614), .S(n5626), .Q(n3274) );
  MUX21X1 U5148 ( .IN1(\R[3][5] ), .IN2(n5615), .S(n5626), .Q(n3273) );
  MUX21X1 U5149 ( .IN1(\R[3][4] ), .IN2(n5616), .S(n5626), .Q(n3272) );
  MUX21X1 U5150 ( .IN1(\R[3][3] ), .IN2(n5617), .S(n5626), .Q(n3271) );
  MUX21X1 U5151 ( .IN1(\R[3][2] ), .IN2(n5618), .S(n5626), .Q(n3270) );
  MUX21X1 U5152 ( .IN1(\R[3][1] ), .IN2(n5619), .S(n5626), .Q(n3269) );
  MUX21X1 U5153 ( .IN1(\R[3][0] ), .IN2(n5620), .S(n5626), .Q(n3268) );
  AND3X1 U5154 ( .IN1(n5621), .IN2(n3806), .IN3(n5717), .Q(n5626) );
  MUX21X1 U5155 ( .IN1(\R[2][31] ), .IN2(n5588), .S(n5627), .Q(n3267) );
  MUX21X1 U5156 ( .IN1(\R[2][30] ), .IN2(n5590), .S(n5627), .Q(n3266) );
  MUX21X1 U5157 ( .IN1(\R[2][29] ), .IN2(n5591), .S(n5627), .Q(n3265) );
  MUX21X1 U5158 ( .IN1(\R[2][28] ), .IN2(n5592), .S(n5627), .Q(n3264) );
  MUX21X1 U5159 ( .IN1(\R[2][27] ), .IN2(n5593), .S(n5627), .Q(n3263) );
  MUX21X1 U5160 ( .IN1(\R[2][26] ), .IN2(n5594), .S(n5627), .Q(n3262) );
  MUX21X1 U5161 ( .IN1(\R[2][25] ), .IN2(n5595), .S(n5627), .Q(n3261) );
  MUX21X1 U5162 ( .IN1(\R[2][24] ), .IN2(n5596), .S(n5627), .Q(n3260) );
  MUX21X1 U5163 ( .IN1(\R[2][23] ), .IN2(n5597), .S(n5627), .Q(n3259) );
  MUX21X1 U5164 ( .IN1(\R[2][22] ), .IN2(n5598), .S(n5627), .Q(n3258) );
  MUX21X1 U5165 ( .IN1(\R[2][21] ), .IN2(n5599), .S(n5627), .Q(n3257) );
  MUX21X1 U5166 ( .IN1(\R[2][20] ), .IN2(n5600), .S(n5627), .Q(n3256) );
  MUX21X1 U5167 ( .IN1(\R[2][19] ), .IN2(n5601), .S(n5627), .Q(n3255) );
  MUX21X1 U5168 ( .IN1(\R[2][18] ), .IN2(n5602), .S(n5627), .Q(n3254) );
  MUX21X1 U5169 ( .IN1(\R[2][17] ), .IN2(n5603), .S(n5627), .Q(n3253) );
  MUX21X1 U5170 ( .IN1(\R[2][16] ), .IN2(n5604), .S(n5627), .Q(n3252) );
  MUX21X1 U5171 ( .IN1(\R[2][15] ), .IN2(n5605), .S(n5627), .Q(n3251) );
  MUX21X1 U5172 ( .IN1(\R[2][14] ), .IN2(n5606), .S(n5627), .Q(n3250) );
  MUX21X1 U5173 ( .IN1(\R[2][13] ), .IN2(n5607), .S(n5627), .Q(n3249) );
  MUX21X1 U5174 ( .IN1(\R[2][12] ), .IN2(n5608), .S(n5627), .Q(n3248) );
  MUX21X1 U5175 ( .IN1(\R[2][11] ), .IN2(n5609), .S(n5627), .Q(n3247) );
  MUX21X1 U5176 ( .IN1(\R[2][10] ), .IN2(n5610), .S(n5627), .Q(n3246) );
  MUX21X1 U5177 ( .IN1(\R[2][9] ), .IN2(n5611), .S(n5627), .Q(n3245) );
  MUX21X1 U5178 ( .IN1(\R[2][8] ), .IN2(n5612), .S(n5627), .Q(n3244) );
  MUX21X1 U5179 ( .IN1(\R[2][7] ), .IN2(n5613), .S(n5627), .Q(n3243) );
  MUX21X1 U5180 ( .IN1(\R[2][6] ), .IN2(n5614), .S(n5627), .Q(n3242) );
  MUX21X1 U5181 ( .IN1(\R[2][5] ), .IN2(n5615), .S(n5627), .Q(n3241) );
  MUX21X1 U5182 ( .IN1(\R[2][4] ), .IN2(n5616), .S(n5627), .Q(n3240) );
  MUX21X1 U5183 ( .IN1(\R[2][3] ), .IN2(n5617), .S(n5627), .Q(n3239) );
  MUX21X1 U5184 ( .IN1(\R[2][2] ), .IN2(n5618), .S(n5627), .Q(n3238) );
  MUX21X1 U5185 ( .IN1(\R[2][1] ), .IN2(n5619), .S(n5627), .Q(n3237) );
  MUX21X1 U5186 ( .IN1(\R[2][0] ), .IN2(n5620), .S(n5627), .Q(n3236) );
  AND3X1 U5187 ( .IN1(n5623), .IN2(n3806), .IN3(n5717), .Q(n5627) );
  MUX21X1 U5188 ( .IN1(\R[1][31] ), .IN2(n5588), .S(n5628), .Q(n3235) );
  MUX21X1 U5189 ( .IN1(\R[1][30] ), .IN2(n5590), .S(n5628), .Q(n3234) );
  MUX21X1 U5190 ( .IN1(\R[1][29] ), .IN2(n5591), .S(n5628), .Q(n3233) );
  MUX21X1 U5191 ( .IN1(\R[1][28] ), .IN2(n5592), .S(n5628), .Q(n3232) );
  MUX21X1 U5192 ( .IN1(\R[1][27] ), .IN2(n5593), .S(n5628), .Q(n3231) );
  MUX21X1 U5193 ( .IN1(\R[1][26] ), .IN2(n5594), .S(n5628), .Q(n3230) );
  MUX21X1 U5194 ( .IN1(\R[1][25] ), .IN2(n5595), .S(n5628), .Q(n3229) );
  MUX21X1 U5195 ( .IN1(\R[1][24] ), .IN2(n5596), .S(n5628), .Q(n3228) );
  MUX21X1 U5196 ( .IN1(\R[1][23] ), .IN2(n5597), .S(n5628), .Q(n3227) );
  MUX21X1 U5197 ( .IN1(\R[1][22] ), .IN2(n5598), .S(n5628), .Q(n3226) );
  MUX21X1 U5198 ( .IN1(\R[1][21] ), .IN2(n5599), .S(n5628), .Q(n3225) );
  MUX21X1 U5199 ( .IN1(\R[1][20] ), .IN2(n5600), .S(n5628), .Q(n3224) );
  MUX21X1 U5200 ( .IN1(\R[1][19] ), .IN2(n5601), .S(n5628), .Q(n3223) );
  MUX21X1 U5201 ( .IN1(\R[1][18] ), .IN2(n5602), .S(n5628), .Q(n3222) );
  MUX21X1 U5202 ( .IN1(\R[1][17] ), .IN2(n5603), .S(n5628), .Q(n3221) );
  MUX21X1 U5203 ( .IN1(\R[1][16] ), .IN2(n5604), .S(n5628), .Q(n3220) );
  MUX21X1 U5204 ( .IN1(\R[1][15] ), .IN2(n5605), .S(n5628), .Q(n3219) );
  MUX21X1 U5205 ( .IN1(\R[1][14] ), .IN2(n5606), .S(n5628), .Q(n3218) );
  MUX21X1 U5206 ( .IN1(\R[1][13] ), .IN2(n5607), .S(n5628), .Q(n3217) );
  MUX21X1 U5207 ( .IN1(\R[1][12] ), .IN2(n5608), .S(n5628), .Q(n3216) );
  MUX21X1 U5208 ( .IN1(\R[1][11] ), .IN2(n5609), .S(n5628), .Q(n3215) );
  MUX21X1 U5209 ( .IN1(\R[1][10] ), .IN2(n5610), .S(n5628), .Q(n3214) );
  MUX21X1 U5210 ( .IN1(\R[1][9] ), .IN2(n5611), .S(n5628), .Q(n3213) );
  MUX21X1 U5211 ( .IN1(\R[1][8] ), .IN2(n5612), .S(n5628), .Q(n3212) );
  MUX21X1 U5212 ( .IN1(\R[1][7] ), .IN2(n5613), .S(n5628), .Q(n3211) );
  MUX21X1 U5213 ( .IN1(\R[1][6] ), .IN2(n5614), .S(n5628), .Q(n3210) );
  MUX21X1 U5214 ( .IN1(\R[1][5] ), .IN2(n5615), .S(n5628), .Q(n3209) );
  MUX21X1 U5215 ( .IN1(\R[1][4] ), .IN2(n5616), .S(n5628), .Q(n3208) );
  MUX21X1 U5216 ( .IN1(\R[1][3] ), .IN2(n5617), .S(n5628), .Q(n3207) );
  MUX21X1 U5217 ( .IN1(\R[1][2] ), .IN2(n5618), .S(n5628), .Q(n3206) );
  MUX21X1 U5218 ( .IN1(\R[1][1] ), .IN2(n5619), .S(n5628), .Q(n3205) );
  MUX21X1 U5219 ( .IN1(\R[1][0] ), .IN2(n5620), .S(n5628), .Q(n3204) );
  AND3X1 U5220 ( .IN1(n5716), .IN2(n5621), .IN3(n5717), .Q(n5628) );
  AND2X1 U5221 ( .IN1(n5629), .IN2(n3883), .Q(n5621) );
  MUX21X1 U5222 ( .IN1(\R[0][31] ), .IN2(n5588), .S(n5630), .Q(n3203) );
  AO22X1 U5223 ( .IN1(n5631), .IN2(n3885), .IN3(data[31]), .IN4(n5632), .Q(
        n5588) );
  MUX21X1 U5224 ( .IN1(\R[0][30] ), .IN2(n5590), .S(n5630), .Q(n3202) );
  AO22X1 U5225 ( .IN1(n5631), .IN2(n3886), .IN3(data[30]), .IN4(n5632), .Q(
        n5590) );
  MUX21X1 U5226 ( .IN1(\R[0][29] ), .IN2(n5591), .S(n5630), .Q(n3201) );
  AO22X1 U5227 ( .IN1(n5631), .IN2(n3887), .IN3(data[29]), .IN4(n5632), .Q(
        n5591) );
  MUX21X1 U5228 ( .IN1(\R[0][28] ), .IN2(n5592), .S(n5630), .Q(n3200) );
  AO22X1 U5229 ( .IN1(n5631), .IN2(n3888), .IN3(data[28]), .IN4(n5632), .Q(
        n5592) );
  MUX21X1 U5230 ( .IN1(\R[0][27] ), .IN2(n5593), .S(n5630), .Q(n3199) );
  AO22X1 U5231 ( .IN1(n5631), .IN2(n3889), .IN3(data[27]), .IN4(n5632), .Q(
        n5593) );
  MUX21X1 U5232 ( .IN1(\R[0][26] ), .IN2(n5594), .S(n5630), .Q(n3198) );
  AO22X1 U5233 ( .IN1(n5631), .IN2(n3890), .IN3(data[26]), .IN4(n5632), .Q(
        n5594) );
  MUX21X1 U5234 ( .IN1(\R[0][25] ), .IN2(n5595), .S(n5630), .Q(n3197) );
  AO22X1 U5235 ( .IN1(n5631), .IN2(n3891), .IN3(data[25]), .IN4(n5632), .Q(
        n5595) );
  MUX21X1 U5236 ( .IN1(\R[0][24] ), .IN2(n5596), .S(n5630), .Q(n3196) );
  AO22X1 U5237 ( .IN1(n5631), .IN2(n3892), .IN3(data[24]), .IN4(n5632), .Q(
        n5596) );
  MUX21X1 U5238 ( .IN1(\R[0][23] ), .IN2(n5597), .S(n5630), .Q(n3195) );
  AO22X1 U5239 ( .IN1(n5631), .IN2(n3893), .IN3(data[23]), .IN4(n5632), .Q(
        n5597) );
  MUX21X1 U5240 ( .IN1(\R[0][22] ), .IN2(n5598), .S(n5630), .Q(n3194) );
  AO22X1 U5241 ( .IN1(n5631), .IN2(n3894), .IN3(data[22]), .IN4(n5632), .Q(
        n5598) );
  MUX21X1 U5242 ( .IN1(\R[0][21] ), .IN2(n5599), .S(n5630), .Q(n3193) );
  AO22X1 U5243 ( .IN1(n5631), .IN2(n3895), .IN3(data[21]), .IN4(n5632), .Q(
        n5599) );
  MUX21X1 U5244 ( .IN1(\R[0][20] ), .IN2(n5600), .S(n5630), .Q(n3192) );
  AO22X1 U5245 ( .IN1(n5631), .IN2(n3896), .IN3(data[20]), .IN4(n5632), .Q(
        n5600) );
  MUX21X1 U5246 ( .IN1(\R[0][19] ), .IN2(n5601), .S(n5630), .Q(n3191) );
  AO22X1 U5247 ( .IN1(n5631), .IN2(n3897), .IN3(data[19]), .IN4(n5632), .Q(
        n5601) );
  MUX21X1 U5248 ( .IN1(\R[0][18] ), .IN2(n5602), .S(n5630), .Q(n3190) );
  AO22X1 U5249 ( .IN1(n5631), .IN2(n3898), .IN3(data[18]), .IN4(n5632), .Q(
        n5602) );
  MUX21X1 U5250 ( .IN1(\R[0][17] ), .IN2(n5603), .S(n5630), .Q(n3189) );
  AO22X1 U5251 ( .IN1(n5631), .IN2(n3899), .IN3(data[17]), .IN4(n5632), .Q(
        n5603) );
  MUX21X1 U5252 ( .IN1(\R[0][16] ), .IN2(n5604), .S(n5630), .Q(n3188) );
  AO22X1 U5253 ( .IN1(n5631), .IN2(n3900), .IN3(data[16]), .IN4(n5632), .Q(
        n5604) );
  MUX21X1 U5254 ( .IN1(\R[0][15] ), .IN2(n5605), .S(n5630), .Q(n3187) );
  AO22X1 U5255 ( .IN1(n5631), .IN2(n3901), .IN3(data[15]), .IN4(n5632), .Q(
        n5605) );
  MUX21X1 U5256 ( .IN1(\R[0][14] ), .IN2(n5606), .S(n5630), .Q(n3186) );
  AO22X1 U5257 ( .IN1(n5631), .IN2(n3902), .IN3(data[14]), .IN4(n5632), .Q(
        n5606) );
  MUX21X1 U5258 ( .IN1(\R[0][13] ), .IN2(n5607), .S(n5630), .Q(n3185) );
  AO22X1 U5259 ( .IN1(n5631), .IN2(n3903), .IN3(data[13]), .IN4(n5632), .Q(
        n5607) );
  MUX21X1 U5260 ( .IN1(\R[0][12] ), .IN2(n5608), .S(n5630), .Q(n3184) );
  AO22X1 U5261 ( .IN1(n5631), .IN2(n3904), .IN3(data[12]), .IN4(n5632), .Q(
        n5608) );
  MUX21X1 U5262 ( .IN1(\R[0][11] ), .IN2(n5609), .S(n5630), .Q(n3183) );
  AO22X1 U5263 ( .IN1(n5631), .IN2(n3905), .IN3(data[11]), .IN4(n5632), .Q(
        n5609) );
  MUX21X1 U5264 ( .IN1(\R[0][10] ), .IN2(n5610), .S(n5630), .Q(n3182) );
  AO22X1 U5265 ( .IN1(n5631), .IN2(n3906), .IN3(data[10]), .IN4(n5632), .Q(
        n5610) );
  MUX21X1 U5266 ( .IN1(\R[0][9] ), .IN2(n5611), .S(n5630), .Q(n3181) );
  AO22X1 U5267 ( .IN1(n5631), .IN2(n3907), .IN3(data[9]), .IN4(n5632), .Q(
        n5611) );
  MUX21X1 U5268 ( .IN1(\R[0][8] ), .IN2(n5612), .S(n5630), .Q(n3180) );
  AO22X1 U5269 ( .IN1(n5631), .IN2(n3908), .IN3(data[8]), .IN4(n5632), .Q(
        n5612) );
  MUX21X1 U5270 ( .IN1(\R[0][7] ), .IN2(n5613), .S(n5630), .Q(n3179) );
  AO22X1 U5271 ( .IN1(n5631), .IN2(n3909), .IN3(data[7]), .IN4(n5632), .Q(
        n5613) );
  MUX21X1 U5272 ( .IN1(\R[0][6] ), .IN2(n5614), .S(n5630), .Q(n3178) );
  AO22X1 U5273 ( .IN1(n5631), .IN2(n3910), .IN3(data[6]), .IN4(n5632), .Q(
        n5614) );
  MUX21X1 U5274 ( .IN1(\R[0][5] ), .IN2(n5615), .S(n5630), .Q(n3177) );
  AO22X1 U5275 ( .IN1(n5631), .IN2(n3911), .IN3(data[5]), .IN4(n5632), .Q(
        n5615) );
  MUX21X1 U5276 ( .IN1(\R[0][4] ), .IN2(n5616), .S(n5630), .Q(n3176) );
  AO22X1 U5277 ( .IN1(n5631), .IN2(n3912), .IN3(data[4]), .IN4(n5632), .Q(
        n5616) );
  MUX21X1 U5278 ( .IN1(\R[0][3] ), .IN2(n5617), .S(n5630), .Q(n3175) );
  AO22X1 U5279 ( .IN1(n5631), .IN2(n3913), .IN3(data[3]), .IN4(n5632), .Q(
        n5617) );
  MUX21X1 U5280 ( .IN1(\R[0][2] ), .IN2(n5618), .S(n5630), .Q(n3174) );
  AO22X1 U5281 ( .IN1(n5631), .IN2(n3914), .IN3(data[2]), .IN4(n5632), .Q(
        n5618) );
  MUX21X1 U5282 ( .IN1(\R[0][1] ), .IN2(n5619), .S(n5630), .Q(n3173) );
  AO22X1 U5283 ( .IN1(n5631), .IN2(n3915), .IN3(data[1]), .IN4(n5632), .Q(
        n5619) );
  MUX21X1 U5284 ( .IN1(\R[0][0] ), .IN2(n5620), .S(n5630), .Q(n3172) );
  AND3X1 U5285 ( .IN1(n5716), .IN2(n5623), .IN3(n5717), .Q(n5630) );
  AND2X1 U5286 ( .IN1(n5714), .IN2(n5629), .Q(n5623) );
  OR2X1 U5287 ( .IN1(n5631), .IN2(n5632), .Q(n5629) );
  AO22X1 U5288 ( .IN1(n5631), .IN2(n3916), .IN3(data[0]), .IN4(n5632), .Q(
        n5620) );
  NOR3X0 U5289 ( .IN1(n5707), .IN2(n5706), .IN3(n5633), .QN(n5632) );
  NAND2X0 U5290 ( .IN1(n5634), .IN2(n5635), .QN(n5631) );
  NAND3X0 U5291 ( .IN1(n5707), .IN2(n5713), .IN3(n5636), .QN(n5635) );
  MUX21X1 U5292 ( .IN1(n5637), .IN2(n5638), .S(n5708), .Q(n5636) );
  NOR3X0 U5293 ( .IN1(n5710), .IN2(n5706), .IN3(n5709), .QN(n5638) );
  INVX0 U5294 ( .INP(n5633), .ZN(n5637) );
  MUX21X1 U5295 ( .IN1(n5639), .IN2(n5640), .S(n5706), .Q(n5634) );
  OA222X1 U5296 ( .IN1(n5641), .IN2(n3846), .IN3(n5642), .IN4(n5643), .IN5(
        n5713), .IN6(n5633), .Q(n5640) );
  NAND2X0 U5297 ( .IN1(n5709), .IN2(n5710), .QN(n5633) );
  OA21X1 U5298 ( .IN1(n5707), .IN2(n5710), .IN3(n3845), .Q(n5642) );
  OA21X1 U5299 ( .IN1(n5644), .IN2(n3882), .IN3(n5645), .Q(n5641) );
  MUX21X1 U5300 ( .IN1(n5646), .IN2(n3884), .S(n5713), .Q(n5645) );
  NAND2X0 U5301 ( .IN1(n5644), .IN2(n3882), .QN(n5646) );
  NOR2X0 U5302 ( .IN1(n5709), .IN2(n5710), .QN(n5644) );
  NAND2X0 U5303 ( .IN1(n5647), .IN2(n3846), .QN(n5639) );
  MUX21X1 U5304 ( .IN1(n5648), .IN2(n5649), .S(n5710), .Q(n5647) );
  AND2X1 U5305 ( .IN1(n3845), .IN2(n5643), .Q(n5649) );
  NAND2X0 U5306 ( .IN1(n5708), .IN2(n5713), .QN(n5643) );
  NOR2X0 U5307 ( .IN1(n5708), .IN2(n3845), .QN(n5648) );
  NOR2X0 U5308 ( .IN1(n5712), .IN2(n5042), .QN(\U3/U76/Z_0 ) );
  NOR2X0 U5309 ( .IN1(n3085), .IN2(n5650), .QN(\U3/U75/Z_9 ) );
  AO22X1 U5310 ( .IN1(n5350), .IN2(ID_imm_offset[6]), .IN3(n5651), .IN4(n4273), 
        .Q(\U3/U75/Z_8 ) );
  INVX0 U5311 ( .INP(n3086), .ZN(n4273) );
  AO222X1 U5312 ( .IN1(n5651), .IN2(n4272), .IN3(n5652), .IN4(ID_imm_offset[7]), .IN5(n5350), .IN6(ID_imm_offset[5]), .Q(\U3/U75/Z_7 ) );
  INVX0 U5313 ( .INP(n3087), .ZN(n4272) );
  AO222X1 U5314 ( .IN1(n5651), .IN2(n4271), .IN3(n5652), .IN4(ID_imm_offset[6]), .IN5(n5350), .IN6(n4371), .Q(\U3/U75/Z_6 ) );
  INVX0 U5315 ( .INP(n3088), .ZN(n4271) );
  AO222X1 U5316 ( .IN1(n5651), .IN2(n4270), .IN3(n5652), .IN4(ID_imm_offset[5]), .IN5(n5350), .IN6(n4375), .Q(\U3/U75/Z_5 ) );
  INVX0 U5317 ( .INP(n3089), .ZN(n4270) );
  AO222X1 U5318 ( .IN1(n5651), .IN2(n4269), .IN3(n5652), .IN4(n4371), .IN5(
        n5350), .IN6(n4381), .Q(\U3/U75/Z_4 ) );
  INVX0 U5319 ( .INP(n2996), .ZN(n4371) );
  INVX0 U5320 ( .INP(n3090), .ZN(n4269) );
  NOR2X0 U5321 ( .IN1(n5725), .IN2(n5650), .QN(\U3/U75/Z_31 ) );
  NOR2X0 U5322 ( .IN1(n3064), .IN2(n5650), .QN(\U3/U75/Z_30 ) );
  AO222X1 U5323 ( .IN1(n5651), .IN2(n4268), .IN3(n5652), .IN4(n4375), .IN5(
        n5350), .IN6(n4383), .Q(\U3/U75/Z_3 ) );
  INVX0 U5324 ( .INP(n2995), .ZN(n4375) );
  INVX0 U5325 ( .INP(n3091), .ZN(n4268) );
  NOR2X0 U5326 ( .IN1(n3065), .IN2(n5650), .QN(\U3/U75/Z_29 ) );
  NOR2X0 U5327 ( .IN1(n3066), .IN2(n5650), .QN(\U3/U75/Z_28 ) );
  NOR2X0 U5328 ( .IN1(n3067), .IN2(n5650), .QN(\U3/U75/Z_27 ) );
  NOR2X0 U5329 ( .IN1(n3068), .IN2(n5650), .QN(\U3/U75/Z_26 ) );
  NOR2X0 U5330 ( .IN1(n3069), .IN2(n5650), .QN(\U3/U75/Z_25 ) );
  NOR2X0 U5331 ( .IN1(n3070), .IN2(n5650), .QN(\U3/U75/Z_24 ) );
  NOR2X0 U5332 ( .IN1(n3071), .IN2(n5650), .QN(\U3/U75/Z_23 ) );
  NOR2X0 U5333 ( .IN1(n3072), .IN2(n5650), .QN(\U3/U75/Z_22 ) );
  NOR2X0 U5334 ( .IN1(n3073), .IN2(n5650), .QN(\U3/U75/Z_21 ) );
  NOR2X0 U5335 ( .IN1(n3074), .IN2(n5650), .QN(\U3/U75/Z_20 ) );
  AO222X1 U5336 ( .IN1(n5651), .IN2(n4267), .IN3(n5653), .IN4(n4381), .IN5(
        n5350), .IN6(n4384), .Q(\U3/U75/Z_2 ) );
  INVX0 U5337 ( .INP(n2994), .ZN(n4381) );
  INVX0 U5338 ( .INP(n3092), .ZN(n4267) );
  NOR2X0 U5339 ( .IN1(n3075), .IN2(n5650), .QN(\U3/U75/Z_19 ) );
  NOR2X0 U5340 ( .IN1(n3076), .IN2(n5650), .QN(\U3/U75/Z_18 ) );
  NOR2X0 U5341 ( .IN1(n3077), .IN2(n5650), .QN(\U3/U75/Z_17 ) );
  NOR2X0 U5342 ( .IN1(n3078), .IN2(n5650), .QN(\U3/U75/Z_16 ) );
  NOR2X0 U5343 ( .IN1(n3079), .IN2(n5650), .QN(\U3/U75/Z_15 ) );
  NOR2X0 U5344 ( .IN1(n3080), .IN2(n5650), .QN(\U3/U75/Z_14 ) );
  NOR2X0 U5345 ( .IN1(n3081), .IN2(n5650), .QN(\U3/U75/Z_13 ) );
  NOR2X0 U5346 ( .IN1(n3082), .IN2(n5650), .QN(\U3/U75/Z_12 ) );
  NOR2X0 U5347 ( .IN1(n3083), .IN2(n5650), .QN(\U3/U75/Z_11 ) );
  NOR2X0 U5348 ( .IN1(n3084), .IN2(n5650), .QN(\U3/U75/Z_10 ) );
  INVX0 U5349 ( .INP(n5651), .ZN(n5650) );
  AO221X1 U5350 ( .IN1(n5653), .IN2(n4383), .IN3(n5651), .IN4(n4266), .IN5(
        n5348), .Q(\U3/U75/Z_1 ) );
  INVX0 U5351 ( .INP(n3093), .ZN(n4266) );
  INVX0 U5352 ( .INP(n2991), .ZN(n4383) );
  AO22X1 U5353 ( .IN1(n5651), .IN2(n4265), .IN3(n5653), .IN4(n4384), .Q(
        \U3/U75/Z_0 ) );
  INVX0 U5354 ( .INP(n2988), .ZN(n4384) );
  NAND2X0 U5355 ( .IN1(n5654), .IN2(n5655), .QN(n5653) );
  INVX0 U5356 ( .INP(n5652), .ZN(n5654) );
  NAND2X0 U5357 ( .IN1(n5074), .IN2(n4582), .QN(n5652) );
  INVX0 U5358 ( .INP(n3094), .ZN(n4265) );
  NAND2X0 U5359 ( .IN1(n5042), .IN2(n5056), .QN(n5651) );
  AO221X1 U5360 ( .IN1(n5656), .IN2(ID_Rn[9]), .IN3(n5657), .IN4(n4335), .IN5(
        n5658), .Q(\U3/U74/Z_9 ) );
  AO22X1 U5361 ( .IN1(n5348), .IN2(ID_PC[9]), .IN3(n5350), .IN4(SP[9]), .Q(
        n5658) );
  INVX0 U5362 ( .INP(n3044), .ZN(n4335) );
  AO221X1 U5363 ( .IN1(n5656), .IN2(ID_Rn[8]), .IN3(n5657), .IN4(n4334), .IN5(
        n5659), .Q(\U3/U74/Z_8 ) );
  AO22X1 U5364 ( .IN1(n5348), .IN2(ID_PC[8]), .IN3(n5350), .IN4(SP[8]), .Q(
        n5659) );
  INVX0 U5365 ( .INP(n3046), .ZN(n4334) );
  AO221X1 U5366 ( .IN1(n5656), .IN2(ID_Rn[7]), .IN3(n5657), .IN4(n4333), .IN5(
        n5660), .Q(\U3/U74/Z_7 ) );
  AO22X1 U5367 ( .IN1(n5348), .IN2(ID_PC[7]), .IN3(n5350), .IN4(SP[7]), .Q(
        n5660) );
  INVX0 U5368 ( .INP(n3048), .ZN(n4333) );
  AO221X1 U5369 ( .IN1(n5656), .IN2(ID_Rn[6]), .IN3(n5657), .IN4(n4332), .IN5(
        n5661), .Q(\U3/U74/Z_6 ) );
  AO22X1 U5370 ( .IN1(n5348), .IN2(ID_PC[6]), .IN3(n5350), .IN4(SP[6]), .Q(
        n5661) );
  INVX0 U5371 ( .INP(n3050), .ZN(n4332) );
  AO221X1 U5372 ( .IN1(n5656), .IN2(ID_Rn[5]), .IN3(n5657), .IN4(n4331), .IN5(
        n5662), .Q(\U3/U74/Z_5 ) );
  AO22X1 U5373 ( .IN1(n5348), .IN2(ID_PC[5]), .IN3(n5350), .IN4(SP[5]), .Q(
        n5662) );
  INVX0 U5374 ( .INP(n3052), .ZN(n4331) );
  AO221X1 U5375 ( .IN1(n5656), .IN2(ID_Rn[4]), .IN3(n5657), .IN4(n4330), .IN5(
        n5663), .Q(\U3/U74/Z_4 ) );
  AO22X1 U5376 ( .IN1(n5348), .IN2(ID_PC[4]), .IN3(n5350), .IN4(SP[4]), .Q(
        n5663) );
  INVX0 U5377 ( .INP(n3054), .ZN(n4330) );
  AO221X1 U5378 ( .IN1(n5656), .IN2(ID_Rn[31]), .IN3(n5657), .IN4(n4357), 
        .IN5(n5664), .Q(\U3/U74/Z_31 ) );
  AO22X1 U5379 ( .IN1(n5348), .IN2(ID_PC[31]), .IN3(n5350), .IN4(SP[31]), .Q(
        n5664) );
  INVX0 U5380 ( .INP(n3000), .ZN(n4357) );
  AO221X1 U5381 ( .IN1(n5656), .IN2(ID_Rn[30]), .IN3(n5657), .IN4(n4356), 
        .IN5(n5665), .Q(\U3/U74/Z_30 ) );
  AO22X1 U5382 ( .IN1(n5348), .IN2(ID_PC[30]), .IN3(n5350), .IN4(SP[30]), .Q(
        n5665) );
  INVX0 U5383 ( .INP(n3002), .ZN(n4356) );
  AO221X1 U5384 ( .IN1(n5656), .IN2(ID_Rn[3]), .IN3(n5657), .IN4(n4329), .IN5(
        n5666), .Q(\U3/U74/Z_3 ) );
  AO22X1 U5385 ( .IN1(n5348), .IN2(ID_PC[3]), .IN3(n5350), .IN4(SP[3]), .Q(
        n5666) );
  INVX0 U5386 ( .INP(n3056), .ZN(n4329) );
  AO221X1 U5387 ( .IN1(n5656), .IN2(ID_Rn[29]), .IN3(n5657), .IN4(n4355), 
        .IN5(n5667), .Q(\U3/U74/Z_29 ) );
  AO22X1 U5388 ( .IN1(n5348), .IN2(ID_PC[29]), .IN3(n5350), .IN4(SP[29]), .Q(
        n5667) );
  INVX0 U5389 ( .INP(n3004), .ZN(n4355) );
  AO221X1 U5390 ( .IN1(n5656), .IN2(ID_Rn[28]), .IN3(n5657), .IN4(n4354), 
        .IN5(n5668), .Q(\U3/U74/Z_28 ) );
  AO22X1 U5391 ( .IN1(n5348), .IN2(ID_PC[28]), .IN3(n5350), .IN4(SP[28]), .Q(
        n5668) );
  INVX0 U5392 ( .INP(n3006), .ZN(n4354) );
  AO221X1 U5393 ( .IN1(n5656), .IN2(ID_Rn[27]), .IN3(n5657), .IN4(n4353), 
        .IN5(n5669), .Q(\U3/U74/Z_27 ) );
  AO22X1 U5394 ( .IN1(n5348), .IN2(ID_PC[27]), .IN3(n5350), .IN4(SP[27]), .Q(
        n5669) );
  INVX0 U5395 ( .INP(n3008), .ZN(n4353) );
  AO221X1 U5396 ( .IN1(n5656), .IN2(ID_Rn[26]), .IN3(n5657), .IN4(n4352), 
        .IN5(n5670), .Q(\U3/U74/Z_26 ) );
  AO22X1 U5397 ( .IN1(n5348), .IN2(ID_PC[26]), .IN3(n5350), .IN4(SP[26]), .Q(
        n5670) );
  INVX0 U5398 ( .INP(n3010), .ZN(n4352) );
  AO221X1 U5399 ( .IN1(n5656), .IN2(ID_Rn[25]), .IN3(n5657), .IN4(n4351), 
        .IN5(n5671), .Q(\U3/U74/Z_25 ) );
  AO22X1 U5400 ( .IN1(n5348), .IN2(ID_PC[25]), .IN3(n5350), .IN4(SP[25]), .Q(
        n5671) );
  INVX0 U5401 ( .INP(n3012), .ZN(n4351) );
  AO221X1 U5402 ( .IN1(n5656), .IN2(ID_Rn[24]), .IN3(n5657), .IN4(n4350), 
        .IN5(n5672), .Q(\U3/U74/Z_24 ) );
  AO22X1 U5403 ( .IN1(n5348), .IN2(ID_PC[24]), .IN3(n5350), .IN4(SP[24]), .Q(
        n5672) );
  INVX0 U5404 ( .INP(n3014), .ZN(n4350) );
  AO221X1 U5405 ( .IN1(n5656), .IN2(ID_Rn[23]), .IN3(n5657), .IN4(n4349), 
        .IN5(n5673), .Q(\U3/U74/Z_23 ) );
  AO22X1 U5406 ( .IN1(n5348), .IN2(ID_PC[23]), .IN3(n5350), .IN4(SP[23]), .Q(
        n5673) );
  INVX0 U5407 ( .INP(n3016), .ZN(n4349) );
  AO221X1 U5408 ( .IN1(n5656), .IN2(ID_Rn[22]), .IN3(n5657), .IN4(n4348), 
        .IN5(n5674), .Q(\U3/U74/Z_22 ) );
  AO22X1 U5409 ( .IN1(n5348), .IN2(ID_PC[22]), .IN3(n5350), .IN4(SP[22]), .Q(
        n5674) );
  INVX0 U5410 ( .INP(n3018), .ZN(n4348) );
  AO221X1 U5411 ( .IN1(n5656), .IN2(ID_Rn[21]), .IN3(n5657), .IN4(n4347), 
        .IN5(n5675), .Q(\U3/U74/Z_21 ) );
  AO22X1 U5412 ( .IN1(n5348), .IN2(ID_PC[21]), .IN3(n5350), .IN4(SP[21]), .Q(
        n5675) );
  INVX0 U5413 ( .INP(n3020), .ZN(n4347) );
  AO221X1 U5414 ( .IN1(n5656), .IN2(ID_Rn[20]), .IN3(n5657), .IN4(n4346), 
        .IN5(n5676), .Q(\U3/U74/Z_20 ) );
  AO22X1 U5415 ( .IN1(n5348), .IN2(ID_PC[20]), .IN3(n5350), .IN4(SP[20]), .Q(
        n5676) );
  INVX0 U5416 ( .INP(n3022), .ZN(n4346) );
  AO221X1 U5417 ( .IN1(n5656), .IN2(ID_Rn[2]), .IN3(n5657), .IN4(n4328), .IN5(
        n5677), .Q(\U3/U74/Z_2 ) );
  AO22X1 U5418 ( .IN1(n5348), .IN2(ID_PC[2]), .IN3(n5350), .IN4(SP[2]), .Q(
        n5677) );
  INVX0 U5419 ( .INP(n3058), .ZN(n4328) );
  AO221X1 U5420 ( .IN1(n5656), .IN2(ID_Rn[19]), .IN3(n5657), .IN4(n4345), 
        .IN5(n5678), .Q(\U3/U74/Z_19 ) );
  AO22X1 U5421 ( .IN1(n5348), .IN2(ID_PC[19]), .IN3(n5350), .IN4(SP[19]), .Q(
        n5678) );
  INVX0 U5422 ( .INP(n3024), .ZN(n4345) );
  AO221X1 U5423 ( .IN1(n5656), .IN2(ID_Rn[18]), .IN3(n5657), .IN4(n4344), 
        .IN5(n5679), .Q(\U3/U74/Z_18 ) );
  AO22X1 U5424 ( .IN1(n5348), .IN2(ID_PC[18]), .IN3(n5350), .IN4(SP[18]), .Q(
        n5679) );
  INVX0 U5425 ( .INP(n3026), .ZN(n4344) );
  AO221X1 U5426 ( .IN1(n5656), .IN2(ID_Rn[17]), .IN3(n5657), .IN4(n4343), 
        .IN5(n5680), .Q(\U3/U74/Z_17 ) );
  AO22X1 U5427 ( .IN1(n5348), .IN2(ID_PC[17]), .IN3(n5350), .IN4(SP[17]), .Q(
        n5680) );
  INVX0 U5428 ( .INP(n3028), .ZN(n4343) );
  AO221X1 U5429 ( .IN1(n5656), .IN2(ID_Rn[16]), .IN3(n5657), .IN4(n4342), 
        .IN5(n5681), .Q(\U3/U74/Z_16 ) );
  AO22X1 U5430 ( .IN1(n5348), .IN2(ID_PC[16]), .IN3(n5350), .IN4(SP[16]), .Q(
        n5681) );
  INVX0 U5431 ( .INP(n3030), .ZN(n4342) );
  AO221X1 U5432 ( .IN1(n5656), .IN2(ID_Rn[15]), .IN3(n5657), .IN4(n4341), 
        .IN5(n5682), .Q(\U3/U74/Z_15 ) );
  AO22X1 U5433 ( .IN1(n5348), .IN2(ID_PC[15]), .IN3(n5350), .IN4(SP[15]), .Q(
        n5682) );
  INVX0 U5434 ( .INP(n3032), .ZN(n4341) );
  AO221X1 U5435 ( .IN1(n5656), .IN2(ID_Rn[14]), .IN3(n5657), .IN4(n4340), 
        .IN5(n5683), .Q(\U3/U74/Z_14 ) );
  AO22X1 U5436 ( .IN1(n5348), .IN2(ID_PC[14]), .IN3(n5350), .IN4(SP[14]), .Q(
        n5683) );
  INVX0 U5437 ( .INP(n3034), .ZN(n4340) );
  AO221X1 U5438 ( .IN1(n5656), .IN2(ID_Rn[13]), .IN3(n5657), .IN4(n4339), 
        .IN5(n5684), .Q(\U3/U74/Z_13 ) );
  AO22X1 U5439 ( .IN1(n5348), .IN2(ID_PC[13]), .IN3(n5350), .IN4(SP[13]), .Q(
        n5684) );
  INVX0 U5440 ( .INP(n3036), .ZN(n4339) );
  AO221X1 U5441 ( .IN1(n5656), .IN2(ID_Rn[12]), .IN3(n5657), .IN4(n4338), 
        .IN5(n5685), .Q(\U3/U74/Z_12 ) );
  AO22X1 U5442 ( .IN1(n5348), .IN2(ID_PC[12]), .IN3(n5350), .IN4(SP[12]), .Q(
        n5685) );
  INVX0 U5443 ( .INP(n3038), .ZN(n4338) );
  AO221X1 U5444 ( .IN1(n5656), .IN2(ID_Rn[11]), .IN3(n5657), .IN4(n4337), 
        .IN5(n5686), .Q(\U3/U74/Z_11 ) );
  AO22X1 U5445 ( .IN1(n5348), .IN2(ID_PC[11]), .IN3(n5350), .IN4(SP[11]), .Q(
        n5686) );
  INVX0 U5446 ( .INP(n3040), .ZN(n4337) );
  AO221X1 U5447 ( .IN1(n5656), .IN2(ID_Rn[10]), .IN3(n5657), .IN4(n4336), 
        .IN5(n5687), .Q(\U3/U74/Z_10 ) );
  AO22X1 U5448 ( .IN1(n5348), .IN2(ID_PC[10]), .IN3(n5350), .IN4(SP[10]), .Q(
        n5687) );
  INVX0 U5449 ( .INP(n3042), .ZN(n4336) );
  AO221X1 U5450 ( .IN1(n5656), .IN2(ID_Rn[1]), .IN3(n5657), .IN4(n4327), .IN5(
        n5688), .Q(\U3/U74/Z_1 ) );
  AO22X1 U5451 ( .IN1(n5348), .IN2(ID_PC[1]), .IN3(n5350), .IN4(SP[1]), .Q(
        n5688) );
  INVX0 U5452 ( .INP(n3060), .ZN(n4327) );
  AO221X1 U5453 ( .IN1(n5656), .IN2(ID_Rn[0]), .IN3(n5657), .IN4(n4325), .IN5(
        n5689), .Q(\U3/U74/Z_0 ) );
  AO22X1 U5454 ( .IN1(n5348), .IN2(ID_PC[0]), .IN3(n5350), .IN4(SP[0]), .Q(
        n5689) );
  NOR2X0 U5455 ( .IN1(n3803), .IN2(n5720), .QN(n5350) );
  INVX0 U5456 ( .INP(n5075), .ZN(n5348) );
  NAND2X0 U5457 ( .IN1(n3807), .IN2(n3803), .QN(n5075) );
  INVX0 U5458 ( .INP(n3062), .ZN(n4325) );
  NAND2X0 U5459 ( .IN1(n4582), .IN2(n5042), .QN(n5657) );
  NAND3X0 U5460 ( .IN1(n5722), .IN2(n5724), .IN3(\r150/A[3] ), .QN(n5042) );
  NAND2X0 U5461 ( .IN1(n5723), .IN2(n3843), .QN(n4582) );
  NAND3X0 U5462 ( .IN1(n5074), .IN2(n5056), .IN3(n5655), .QN(n5656) );
  OA22X1 U5463 ( .IN1(n3804), .IN2(\r150/A[3] ), .IN3(n3843), .IN4(n5723), .Q(
        n5655) );
  NAND2X0 U5464 ( .IN1(n3843), .IN2(n3803), .QN(n5056) );
  NAND2X0 U5465 ( .IN1(\r150/A[3] ), .IN2(n3805), .QN(n5074) );
  NAND2X0 U5466 ( .IN1(N695), .IN2(N694), .QN(N693) );
  NAND2X0 U5467 ( .IN1(n5719), .IN2(n5690), .QN(N694) );
  NAND2X0 U5468 ( .IN1(n5690), .IN2(n4369), .QN(N695) );
  NOR3X0 U5469 ( .IN1(n5727), .IN2(n5726), .IN3(n3799), .QN(n5690) );
  AO21X1 U5470 ( .IN1(n4368), .IN2(n4369), .IN3(n3797), .Q(N690) );
  OA21X1 U5471 ( .IN1(n4260), .IN2(n5691), .IN3(n5692), .Q(N688) );
  OAI21X1 U5472 ( .IN1(n4245), .IN2(n5693), .IN3(IF_IR[12]), .QN(N687) );
  NOR2X0 U5473 ( .IN1(n5737), .IN2(n5693), .QN(N686) );
  AO21X1 U5474 ( .IN1(n5691), .IN2(n5692), .IN3(n3802), .Q(N685) );
  NAND3X0 U5475 ( .IN1(n4306), .IN2(n5694), .IN3(n5695), .QN(N599) );
  NAND2X0 U5476 ( .IN1(n4320), .IN2(n5739), .QN(n5695) );
  INVX0 U5477 ( .INP(n4389), .ZN(n4320) );
  OR2X1 U5478 ( .IN1(n4368), .IN2(N598), .Q(N596) );
  NAND3X0 U5479 ( .IN1(n4319), .IN2(n4304), .IN3(n4389), .QN(N598) );
  INVX0 U5480 ( .INP(n4306), .ZN(n4368) );
  NAND3X0 U5481 ( .IN1(n4319), .IN2(n4306), .IN3(n4389), .QN(N595) );
  NAND3X0 U5482 ( .IN1(n4306), .IN2(n4304), .IN3(n4299), .QN(n4389) );
  AND3X1 U5483 ( .IN1(n4319), .IN2(n5694), .IN3(n4318), .Q(n4299) );
  NAND4X0 U5484 ( .IN1(n5696), .IN2(n5697), .IN3(n5719), .IN4(n5698), .QN(
        n4318) );
  NOR2X0 U5485 ( .IN1(n5699), .IN2(n4260), .QN(n5698) );
  INVX0 U5486 ( .INP(n3096), .ZN(n4260) );
  NAND3X0 U5487 ( .IN1(n5693), .IN2(n5705), .IN3(n5700), .QN(n5694) );
  OR2X1 U5488 ( .IN1(n4241), .IN2(n3795), .Q(n4304) );
  NAND2X0 U5489 ( .IN1(n5696), .IN2(n5692), .QN(n4306) );
  INVX0 U5490 ( .INP(n5737), .ZN(n5692) );
  NAND2X0 U5491 ( .IN1(n3799), .IN2(IF_IR[12]), .QN(n5737) );
  NAND3X0 U5492 ( .IN1(n5693), .IN2(n5697), .IN3(n5700), .QN(n4319) );
  INVX0 U5493 ( .INP(n5705), .ZN(n5697) );
  NOR2X0 U5494 ( .IN1(n5691), .IN2(n3096), .QN(n5693) );
  NAND2X0 U5495 ( .IN1(n5696), .IN2(n4369), .QN(n5691) );
  INVX0 U5496 ( .INP(n5719), .ZN(n4369) );
  NOR2X0 U5497 ( .IN1(n4241), .IN2(n4243), .QN(n5696) );
  INVX0 U5498 ( .INP(n5726), .ZN(n4243) );
  AO21X1 U5499 ( .IN1(n4245), .IN2(n4241), .IN3(n3802), .Q(N550) );
  INVX0 U5500 ( .INP(n5739), .ZN(n3802) );
  NAND2X0 U5501 ( .IN1(n3797), .IN2(n4245), .QN(n5739) );
  AO21X1 U5502 ( .IN1(N498), .IN2(n4241), .IN3(n5700), .Q(N548) );
  INVX0 U5503 ( .INP(n5699), .ZN(n5700) );
  INVX0 U5504 ( .INP(n5727), .ZN(n4241) );
  NAND2X0 U5505 ( .IN1(n3795), .IN2(n5699), .QN(N547) );
  NAND2X0 U5506 ( .IN1(n3797), .IN2(n3799), .QN(n5699) );
  NAND2X0 U5507 ( .IN1(n5726), .IN2(N498), .QN(n3795) );
  INVX0 U5508 ( .INP(n5738), .ZN(N498) );
  NAND2X0 U5509 ( .IN1(IF_IR[12]), .IN2(n4245), .QN(n5738) );
  INVX0 U5510 ( .INP(n3799), .ZN(n4245) );
  NAND3X0 U5511 ( .IN1(n5721), .IN2(n5711), .IN3(n5701), .QN(N4637) );
  OA221X1 U5512 ( .IN1(n3805), .IN2(n3807), .IN3(n4406), .IN4(n5073), .IN5(
        n3804), .Q(n5701) );
  INVX0 U5513 ( .INP(n4429), .ZN(n4406) );
  NAND2X0 U5514 ( .IN1(n5721), .IN2(n5720), .QN(n4429) );
  NAND4X0 U5515 ( .IN1(n5702), .IN2(n5711), .IN3(n5703), .IN4(n3844), .QN(
        N4634) );
  NAND2X0 U5516 ( .IN1(n5704), .IN2(n5073), .QN(n5703) );
  AO21X1 U5517 ( .IN1(n3805), .IN2(n3803), .IN3(n3807), .Q(n5704) );
  MUX21X1 U5518 ( .IN1(n5073), .IN2(n3807), .S(n5722), .Q(n5702) );
  NAND2X0 U5519 ( .IN1(n3843), .IN2(n3805), .QN(n5073) );
  MUX21X1 U5520 ( .IN1(N232), .IN2(n3848), .S(n3842), .Q(N344) );
  MUX21X1 U5521 ( .IN1(N231), .IN2(n3849), .S(n3842), .Q(N343) );
  MUX21X1 U5522 ( .IN1(N230), .IN2(n3850), .S(n3842), .Q(N342) );
  MUX21X1 U5523 ( .IN1(N229), .IN2(n3851), .S(n3842), .Q(N341) );
  MUX21X1 U5524 ( .IN1(N228), .IN2(n3852), .S(n3842), .Q(N340) );
  MUX21X1 U5525 ( .IN1(N227), .IN2(n3853), .S(n3842), .Q(N339) );
  MUX21X1 U5526 ( .IN1(N226), .IN2(n3854), .S(n3842), .Q(N338) );
  MUX21X1 U5527 ( .IN1(N225), .IN2(n3855), .S(n3842), .Q(N337) );
  MUX21X1 U5528 ( .IN1(N224), .IN2(n3856), .S(n3842), .Q(N336) );
  MUX21X1 U5529 ( .IN1(N223), .IN2(n3857), .S(n3842), .Q(N335) );
  MUX21X1 U5530 ( .IN1(N222), .IN2(n3858), .S(n3842), .Q(N334) );
  MUX21X1 U5531 ( .IN1(N221), .IN2(n3859), .S(n3842), .Q(N333) );
  MUX21X1 U5532 ( .IN1(N220), .IN2(n3860), .S(n3842), .Q(N332) );
  MUX21X1 U5533 ( .IN1(N219), .IN2(n3861), .S(n3842), .Q(N331) );
  MUX21X1 U5534 ( .IN1(N218), .IN2(n3862), .S(n3842), .Q(N330) );
  MUX21X1 U5535 ( .IN1(N217), .IN2(n3863), .S(n3842), .Q(N329) );
  MUX21X1 U5536 ( .IN1(N216), .IN2(n3864), .S(n3842), .Q(N328) );
  MUX21X1 U5537 ( .IN1(N215), .IN2(n3865), .S(n3842), .Q(N327) );
  MUX21X1 U5538 ( .IN1(N214), .IN2(n3866), .S(n3842), .Q(N326) );
  MUX21X1 U5539 ( .IN1(N213), .IN2(n3867), .S(n3842), .Q(N325) );
  MUX21X1 U5540 ( .IN1(N212), .IN2(n3868), .S(n3842), .Q(N324) );
  MUX21X1 U5541 ( .IN1(N211), .IN2(n3869), .S(n3842), .Q(N323) );
  MUX21X1 U5542 ( .IN1(N210), .IN2(n3870), .S(n3842), .Q(N322) );
  MUX21X1 U5543 ( .IN1(N209), .IN2(n3871), .S(n3842), .Q(N321) );
  MUX21X1 U5544 ( .IN1(N208), .IN2(n3872), .S(n3842), .Q(N320) );
  MUX21X1 U5545 ( .IN1(N207), .IN2(n3873), .S(n3842), .Q(N319) );
  MUX21X1 U5546 ( .IN1(N206), .IN2(n3874), .S(n3842), .Q(N318) );
  MUX21X1 U5547 ( .IN1(N205), .IN2(n3875), .S(n3842), .Q(N317) );
  MUX21X1 U5548 ( .IN1(N204), .IN2(n3876), .S(n3842), .Q(N316) );
  MUX21X1 U5549 ( .IN1(N203), .IN2(n3877), .S(n3842), .Q(N315) );
  MUX21X1 U5550 ( .IN1(N202), .IN2(n3878), .S(n3842), .Q(N314) );
  MUX21X1 U5551 ( .IN1(N201), .IN2(n3879), .S(n3842), .Q(N313) );
endmodule


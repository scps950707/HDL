
module pipealu_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403;

  INVX0 U655 ( .INP(n1337), .ZN(n1296) );
  INVX0 U656 ( .INP(n1373), .ZN(n1280) );
  INVX0 U657 ( .INP(n1327), .ZN(n1288) );
  INVX0 U658 ( .INP(n1372), .ZN(n1285) );
  INVX0 U659 ( .INP(n1371), .ZN(n1281) );
  INVX0 U660 ( .INP(n1332), .ZN(n1294) );
  INVX0 U661 ( .INP(n1394), .ZN(n1290) );
  INVX0 U662 ( .INP(B[20]), .ZN(n1291) );
  INVX0 U663 ( .INP(n1347), .ZN(n1297) );
  INVX0 U664 ( .INP(n1383), .ZN(n1282) );
  INVX0 U665 ( .INP(n1338), .ZN(n1300) );
  OR3X1 U666 ( .IN1(n1358), .IN2(n1278), .IN3(n1279), .Q(n1339) );
  AOI221X1 U667 ( .IN1(B[1]), .IN2(n1321), .IN3(n1366), .IN4(B[0]), .IN5(n1364), .QN(n1278) );
  OAI221X1 U668 ( .IN1(n1363), .IN2(n1364), .IN3(B[4]), .IN4(n1319), .IN5(
        n1362), .QN(n1279) );
  INVX0 U669 ( .INP(B[18]), .ZN(n1293) );
  INVX0 U670 ( .INP(A[12]), .ZN(n1315) );
  INVX0 U671 ( .INP(A[8]), .ZN(n1317) );
  INVX0 U672 ( .INP(A[28]), .ZN(n1307) );
  INVX0 U673 ( .INP(A[24]), .ZN(n1309) );
  INVX0 U674 ( .INP(A[31]), .ZN(n1306) );
  INVX0 U675 ( .INP(B[14]), .ZN(n1298) );
  INVX0 U676 ( .INP(B[6]), .ZN(n1303) );
  INVX0 U677 ( .INP(B[30]), .ZN(n1283) );
  INVX0 U678 ( .INP(B[10]), .ZN(n1301) );
  INVX0 U679 ( .INP(B[26]), .ZN(n1286) );
  INVX0 U680 ( .INP(A[4]), .ZN(n1319) );
  INVX0 U681 ( .INP(A[21]), .ZN(n1311) );
  INVX0 U682 ( .INP(A[17]), .ZN(n1313) );
  INVX0 U683 ( .INP(A[3]), .ZN(n1320) );
  INVX0 U684 ( .INP(A[23]), .ZN(n1310) );
  INVX0 U685 ( .INP(A[19]), .ZN(n1312) );
  INVX0 U686 ( .INP(A[1]), .ZN(n1321) );
  INVX0 U687 ( .INP(A[11]), .ZN(n1316) );
  INVX0 U688 ( .INP(A[15]), .ZN(n1314) );
  INVX0 U689 ( .INP(A[27]), .ZN(n1308) );
  INVX0 U690 ( .INP(A[7]), .ZN(n1318) );
  INVX0 U691 ( .INP(B[9]), .ZN(n1302) );
  INVX0 U692 ( .INP(B[13]), .ZN(n1299) );
  INVX0 U693 ( .INP(B[5]), .ZN(n1304) );
  INVX0 U694 ( .INP(B[25]), .ZN(n1287) );
  INVX0 U695 ( .INP(B[29]), .ZN(n1284) );
  INVX0 U696 ( .INP(n1326), .ZN(n1292) );
  INVX0 U697 ( .INP(B[22]), .ZN(n1289) );
  INVX0 U698 ( .INP(B[2]), .ZN(n1305) );
  INVX0 U699 ( .INP(B[16]), .ZN(n1295) );
  AO21X1 U700 ( .IN1(n1322), .IN2(n1323), .IN3(n1324), .Q(GE_LT_GT_LE) );
  NOR4X0 U701 ( .IN1(n1325), .IN2(n1326), .IN3(n1327), .IN4(n1328), .QN(n1324)
         );
  NAND4X0 U702 ( .IN1(n1329), .IN2(n1330), .IN3(n1294), .IN4(n1331), .QN(n1325) );
  NAND2X0 U703 ( .IN1(A[16]), .IN2(n1295), .QN(n1331) );
  NAND2X0 U704 ( .IN1(n1333), .IN2(n1334), .QN(n1330) );
  NAND4X0 U705 ( .IN1(n1300), .IN2(n1296), .IN3(n1335), .IN4(n1336), .QN(n1334) );
  OR2X1 U706 ( .IN1(n1317), .IN2(B[8]), .Q(n1336) );
  NAND3X0 U707 ( .IN1(n1339), .IN2(n1340), .IN3(n1333), .QN(n1329) );
  AND2X1 U708 ( .IN1(n1341), .IN2(n1342), .Q(n1333) );
  AO221X1 U709 ( .IN1(n1343), .IN2(n1338), .IN3(n1344), .IN4(n1343), .IN5(
        n1337), .Q(n1342) );
  NAND3X0 U710 ( .IN1(n1345), .IN2(n1346), .IN3(n1297), .QN(n1337) );
  OR2X1 U711 ( .IN1(n1315), .IN2(B[12]), .Q(n1346) );
  OA21X1 U712 ( .IN1(A[9]), .IN2(n1302), .IN3(n1348), .Q(n1344) );
  NAND3X0 U713 ( .IN1(n1335), .IN2(n1317), .IN3(B[8]), .QN(n1348) );
  NAND2X0 U714 ( .IN1(A[9]), .IN2(n1302), .QN(n1335) );
  AO21X1 U715 ( .IN1(A[10]), .IN2(n1301), .IN3(n1349), .Q(n1338) );
  AOI22X1 U716 ( .IN1(B[11]), .IN2(n1316), .IN3(n1350), .IN4(B[10]), .QN(n1343) );
  NOR2X0 U717 ( .IN1(A[10]), .IN2(n1349), .QN(n1350) );
  NOR2X0 U718 ( .IN1(n1316), .IN2(B[11]), .QN(n1349) );
  AO22X1 U719 ( .IN1(n1351), .IN2(n1352), .IN3(n1352), .IN4(n1347), .Q(n1341)
         );
  AO21X1 U720 ( .IN1(A[14]), .IN2(n1298), .IN3(n1353), .Q(n1347) );
  AOI22X1 U721 ( .IN1(B[15]), .IN2(n1314), .IN3(n1354), .IN4(B[14]), .QN(n1352) );
  NOR2X0 U722 ( .IN1(A[14]), .IN2(n1353), .QN(n1354) );
  NOR2X0 U723 ( .IN1(n1314), .IN2(B[15]), .QN(n1353) );
  OA21X1 U724 ( .IN1(A[13]), .IN2(n1299), .IN3(n1355), .Q(n1351) );
  NAND3X0 U725 ( .IN1(n1345), .IN2(n1315), .IN3(B[12]), .QN(n1355) );
  NAND2X0 U726 ( .IN1(A[13]), .IN2(n1299), .QN(n1345) );
  AO22X1 U727 ( .IN1(n1356), .IN2(n1357), .IN3(n1357), .IN4(n1358), .Q(n1340)
         );
  AOI22X1 U728 ( .IN1(B[7]), .IN2(n1318), .IN3(n1359), .IN4(B[6]), .QN(n1357)
         );
  NOR2X0 U729 ( .IN1(A[6]), .IN2(n1360), .QN(n1359) );
  OA21X1 U730 ( .IN1(A[5]), .IN2(n1304), .IN3(n1361), .Q(n1356) );
  NAND3X0 U731 ( .IN1(n1362), .IN2(n1319), .IN3(B[4]), .QN(n1361) );
  NAND2X0 U732 ( .IN1(A[5]), .IN2(n1304), .QN(n1362) );
  AOI21X1 U733 ( .IN1(n1305), .IN2(A[2]), .IN3(n1365), .QN(n1363) );
  AO22X1 U734 ( .IN1(B[3]), .IN2(n1320), .IN3(n1367), .IN4(B[2]), .Q(n1364) );
  NOR2X0 U735 ( .IN1(A[2]), .IN2(n1365), .QN(n1367) );
  NOR2X0 U736 ( .IN1(n1320), .IN2(B[3]), .QN(n1365) );
  NOR2X0 U737 ( .IN1(A[0]), .IN2(n1368), .QN(n1366) );
  NOR2X0 U738 ( .IN1(B[1]), .IN2(n1321), .QN(n1368) );
  AO21X1 U739 ( .IN1(A[6]), .IN2(n1303), .IN3(n1360), .Q(n1358) );
  NOR2X0 U740 ( .IN1(n1318), .IN2(B[7]), .QN(n1360) );
  NAND2X0 U741 ( .IN1(n1280), .IN2(n1328), .QN(n1323) );
  NAND4X0 U742 ( .IN1(n1285), .IN2(n1281), .IN3(n1369), .IN4(n1370), .QN(n1328) );
  OR2X1 U743 ( .IN1(n1309), .IN2(B[24]), .Q(n1370) );
  AO221X1 U744 ( .IN1(n1374), .IN2(n1375), .IN3(n1376), .IN4(n1288), .IN5(
        n1373), .Q(n1322) );
  NAND2X0 U745 ( .IN1(n1377), .IN2(n1378), .QN(n1373) );
  AO221X1 U746 ( .IN1(n1379), .IN2(n1372), .IN3(n1380), .IN4(n1379), .IN5(
        n1371), .Q(n1378) );
  NAND3X0 U747 ( .IN1(n1381), .IN2(n1382), .IN3(n1282), .QN(n1371) );
  OR2X1 U748 ( .IN1(n1307), .IN2(B[28]), .Q(n1382) );
  OA21X1 U749 ( .IN1(A[25]), .IN2(n1287), .IN3(n1384), .Q(n1380) );
  NAND3X0 U750 ( .IN1(n1369), .IN2(n1309), .IN3(B[24]), .QN(n1384) );
  NAND2X0 U751 ( .IN1(A[25]), .IN2(n1287), .QN(n1369) );
  AO21X1 U752 ( .IN1(A[26]), .IN2(n1286), .IN3(n1385), .Q(n1372) );
  AOI22X1 U753 ( .IN1(B[27]), .IN2(n1308), .IN3(n1386), .IN4(B[26]), .QN(n1379) );
  NOR2X0 U754 ( .IN1(A[26]), .IN2(n1385), .QN(n1386) );
  NOR2X0 U755 ( .IN1(n1308), .IN2(B[27]), .QN(n1385) );
  AO22X1 U756 ( .IN1(n1387), .IN2(n1388), .IN3(n1388), .IN4(n1383), .Q(n1377)
         );
  AO21X1 U757 ( .IN1(A[30]), .IN2(n1283), .IN3(n1389), .Q(n1383) );
  AOI22X1 U758 ( .IN1(B[31]), .IN2(n1306), .IN3(n1390), .IN4(B[30]), .QN(n1388) );
  NOR2X0 U759 ( .IN1(A[30]), .IN2(n1389), .QN(n1390) );
  NOR2X0 U760 ( .IN1(n1306), .IN2(B[31]), .QN(n1389) );
  OA21X1 U761 ( .IN1(A[29]), .IN2(n1284), .IN3(n1391), .Q(n1387) );
  NAND3X0 U762 ( .IN1(n1381), .IN2(n1307), .IN3(B[28]), .QN(n1391) );
  NAND2X0 U763 ( .IN1(A[29]), .IN2(n1284), .QN(n1381) );
  NAND3X0 U764 ( .IN1(n1290), .IN2(n1392), .IN3(n1393), .QN(n1327) );
  NAND2X0 U765 ( .IN1(A[20]), .IN2(n1291), .QN(n1392) );
  OA21X1 U766 ( .IN1(n1292), .IN2(n1395), .IN3(n1396), .Q(n1376) );
  AO221X1 U767 ( .IN1(B[17]), .IN2(n1313), .IN3(n1397), .IN4(B[16]), .IN5(
        n1395), .Q(n1396) );
  NOR2X0 U768 ( .IN1(A[16]), .IN2(n1332), .QN(n1397) );
  NOR2X0 U769 ( .IN1(n1313), .IN2(B[17]), .QN(n1332) );
  AO22X1 U770 ( .IN1(B[19]), .IN2(n1312), .IN3(n1398), .IN4(B[18]), .Q(n1395)
         );
  NOR2X0 U771 ( .IN1(A[18]), .IN2(n1399), .QN(n1398) );
  AO21X1 U772 ( .IN1(A[18]), .IN2(n1293), .IN3(n1399), .Q(n1326) );
  NOR2X0 U773 ( .IN1(n1312), .IN2(B[19]), .QN(n1399) );
  OR2X1 U774 ( .IN1(n1400), .IN2(n1393), .Q(n1375) );
  AOI21X1 U775 ( .IN1(A[22]), .IN2(n1289), .IN3(n1401), .QN(n1393) );
  AO221X1 U776 ( .IN1(B[21]), .IN2(n1311), .IN3(n1402), .IN4(B[20]), .IN5(
        n1400), .Q(n1374) );
  AO22X1 U777 ( .IN1(B[23]), .IN2(n1310), .IN3(n1403), .IN4(B[22]), .Q(n1400)
         );
  NOR2X0 U778 ( .IN1(A[22]), .IN2(n1401), .QN(n1403) );
  NOR2X0 U779 ( .IN1(n1310), .IN2(B[23]), .QN(n1401) );
  NOR2X0 U780 ( .IN1(A[20]), .IN2(n1394), .QN(n1402) );
  NOR2X0 U781 ( .IN1(n1311), .IN2(B[21]), .QN(n1394) );
endmodule


module pipealu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;
  wire   [33:0] carry;

  FADDX1 U2_31 ( .A(A[31]), .B(n4), .CI(carry[31]), .CO(carry[32]), .S(
        DIFF[31]) );
  FADDX1 U2_30 ( .A(A[30]), .B(n5), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  FADDX1 U2_29 ( .A(A[29]), .B(n6), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  FADDX1 U2_28 ( .A(A[28]), .B(n7), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  FADDX1 U2_27 ( .A(A[27]), .B(n8), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  FADDX1 U2_26 ( .A(A[26]), .B(n9), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  FADDX1 U2_25 ( .A(A[25]), .B(n10), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  FADDX1 U2_24 ( .A(A[24]), .B(n11), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  FADDX1 U2_23 ( .A(A[23]), .B(n12), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1 U2_22 ( .A(A[22]), .B(n13), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n14), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n15), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n16), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n17), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n18), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n19), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n20), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n21), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n22), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n23), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n24), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n25), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n26), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n27), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_7 ( .A(A[7]), .B(n28), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  FADDX1 U2_6 ( .A(A[6]), .B(n29), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FADDX1 U2_5 ( .A(A[5]), .B(n30), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  FADDX1 U2_4 ( .A(A[4]), .B(n31), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  FADDX1 U2_3 ( .A(A[3]), .B(n32), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n33), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n34), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  INVX0 U1 ( .INP(carry[32]), .ZN(DIFF[32]) );
  INVX0 U2 ( .INP(B[6]), .ZN(n29) );
  INVX0 U3 ( .INP(B[10]), .ZN(n25) );
  INVX0 U4 ( .INP(B[14]), .ZN(n21) );
  INVX0 U5 ( .INP(B[18]), .ZN(n17) );
  INVX0 U6 ( .INP(B[26]), .ZN(n9) );
  INVX0 U7 ( .INP(B[30]), .ZN(n5) );
  INVX0 U8 ( .INP(B[16]), .ZN(n19) );
  INVX0 U9 ( .INP(B[20]), .ZN(n15) );
  INVX0 U10 ( .INP(B[22]), .ZN(n13) );
  INVX0 U11 ( .INP(B[2]), .ZN(n33) );
  INVX0 U12 ( .INP(B[1]), .ZN(n34) );
  NAND2X1 U13 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U14 ( .INP(A[0]), .ZN(n1) );
  INVX0 U15 ( .INP(B[3]), .ZN(n32) );
  INVX0 U16 ( .INP(B[4]), .ZN(n31) );
  INVX0 U17 ( .INP(B[7]), .ZN(n28) );
  INVX0 U18 ( .INP(B[8]), .ZN(n27) );
  INVX0 U19 ( .INP(B[11]), .ZN(n24) );
  INVX0 U20 ( .INP(B[12]), .ZN(n23) );
  INVX0 U21 ( .INP(B[15]), .ZN(n20) );
  INVX0 U22 ( .INP(B[17]), .ZN(n18) );
  INVX0 U23 ( .INP(B[19]), .ZN(n16) );
  INVX0 U24 ( .INP(B[21]), .ZN(n14) );
  INVX0 U25 ( .INP(B[23]), .ZN(n12) );
  INVX0 U26 ( .INP(B[24]), .ZN(n11) );
  INVX0 U27 ( .INP(B[27]), .ZN(n8) );
  INVX0 U28 ( .INP(B[28]), .ZN(n7) );
  INVX0 U29 ( .INP(B[5]), .ZN(n30) );
  INVX0 U30 ( .INP(B[13]), .ZN(n22) );
  INVX0 U31 ( .INP(B[25]), .ZN(n10) );
  INVX0 U32 ( .INP(B[29]), .ZN(n6) );
  INVX0 U33 ( .INP(B[9]), .ZN(n26) );
  INVX0 U34 ( .INP(B[31]), .ZN(n4) );
  INVX0 U35 ( .INP(n35), .ZN(n2) );
  INVX0 U36 ( .INP(B[0]), .ZN(n35) );
  XOR2X1 U37 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module pipealu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [32:1] carry;

  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(SUM[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module pipealu ( instr, AluOut, Zero, clk, Carryout, Overflow );
  input [15:0] instr;
  output [31:0] AluOut;
  input clk;
  output Zero, Carryout, Overflow;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, \regfile[15][31] ,
         \regfile[15][30] , \regfile[15][29] , \regfile[15][28] ,
         \regfile[15][27] , \regfile[15][26] , \regfile[15][25] ,
         \regfile[15][24] , \regfile[15][23] , \regfile[15][22] ,
         \regfile[15][21] , \regfile[15][20] , \regfile[15][19] ,
         \regfile[15][18] , \regfile[15][17] , \regfile[15][16] ,
         \regfile[15][15] , \regfile[15][14] , \regfile[15][13] ,
         \regfile[15][12] , \regfile[15][11] , \regfile[15][10] ,
         \regfile[15][9] , \regfile[15][8] , \regfile[15][7] ,
         \regfile[15][6] , \regfile[15][5] , \regfile[15][4] ,
         \regfile[15][3] , \regfile[15][2] , \regfile[15][1] ,
         \regfile[15][0] , \regfile[14][31] , \regfile[14][30] ,
         \regfile[14][29] , \regfile[14][28] , \regfile[14][27] ,
         \regfile[14][26] , \regfile[14][25] , \regfile[14][24] ,
         \regfile[14][23] , \regfile[14][22] , \regfile[14][21] ,
         \regfile[14][20] , \regfile[14][19] , \regfile[14][18] ,
         \regfile[14][17] , \regfile[14][16] , \regfile[14][15] ,
         \regfile[14][14] , \regfile[14][13] , \regfile[14][12] ,
         \regfile[14][11] , \regfile[14][10] , \regfile[14][9] ,
         \regfile[14][8] , \regfile[14][7] , \regfile[14][6] ,
         \regfile[14][5] , \regfile[14][4] , \regfile[14][3] ,
         \regfile[14][2] , \regfile[14][1] , \regfile[14][0] ,
         \regfile[13][31] , \regfile[13][30] , \regfile[13][29] ,
         \regfile[13][28] , \regfile[13][27] , \regfile[13][26] ,
         \regfile[13][25] , \regfile[13][24] , \regfile[13][23] ,
         \regfile[13][22] , \regfile[13][21] , \regfile[13][20] ,
         \regfile[13][19] , \regfile[13][18] , \regfile[13][17] ,
         \regfile[13][16] , \regfile[13][15] , \regfile[13][14] ,
         \regfile[13][13] , \regfile[13][12] , \regfile[13][11] ,
         \regfile[13][10] , \regfile[13][9] , \regfile[13][8] ,
         \regfile[13][7] , \regfile[13][6] , \regfile[13][5] ,
         \regfile[13][4] , \regfile[13][3] , \regfile[13][2] ,
         \regfile[13][1] , \regfile[13][0] , \regfile[12][31] ,
         \regfile[12][30] , \regfile[12][29] , \regfile[12][28] ,
         \regfile[12][27] , \regfile[12][26] , \regfile[12][25] ,
         \regfile[12][24] , \regfile[12][23] , \regfile[12][22] ,
         \regfile[12][21] , \regfile[12][20] , \regfile[12][19] ,
         \regfile[12][18] , \regfile[12][17] , \regfile[12][16] ,
         \regfile[12][15] , \regfile[12][14] , \regfile[12][13] ,
         \regfile[12][12] , \regfile[12][11] , \regfile[12][10] ,
         \regfile[12][9] , \regfile[12][8] , \regfile[12][7] ,
         \regfile[12][6] , \regfile[12][5] , \regfile[12][4] ,
         \regfile[12][3] , \regfile[12][2] , \regfile[12][1] ,
         \regfile[12][0] , \regfile[11][31] , \regfile[11][30] ,
         \regfile[11][29] , \regfile[11][28] , \regfile[11][27] ,
         \regfile[11][26] , \regfile[11][25] , \regfile[11][24] ,
         \regfile[11][23] , \regfile[11][22] , \regfile[11][21] ,
         \regfile[11][20] , \regfile[11][19] , \regfile[11][18] ,
         \regfile[11][17] , \regfile[11][16] , \regfile[11][15] ,
         \regfile[11][14] , \regfile[11][13] , \regfile[11][12] ,
         \regfile[11][11] , \regfile[11][10] , \regfile[11][9] ,
         \regfile[11][8] , \regfile[11][7] , \regfile[11][6] ,
         \regfile[11][5] , \regfile[11][4] , \regfile[11][3] ,
         \regfile[11][2] , \regfile[11][1] , \regfile[11][0] ,
         \regfile[10][31] , \regfile[10][30] , \regfile[10][29] ,
         \regfile[10][28] , \regfile[10][27] , \regfile[10][26] ,
         \regfile[10][25] , \regfile[10][24] , \regfile[10][23] ,
         \regfile[10][22] , \regfile[10][21] , \regfile[10][20] ,
         \regfile[10][19] , \regfile[10][18] , \regfile[10][17] ,
         \regfile[10][16] , \regfile[10][15] , \regfile[10][14] ,
         \regfile[10][13] , \regfile[10][12] , \regfile[10][11] ,
         \regfile[10][10] , \regfile[10][9] , \regfile[10][8] ,
         \regfile[10][7] , \regfile[10][6] , \regfile[10][5] ,
         \regfile[10][4] , \regfile[10][3] , \regfile[10][2] ,
         \regfile[10][1] , \regfile[10][0] , \regfile[9][31] ,
         \regfile[9][30] , \regfile[9][29] , \regfile[9][28] ,
         \regfile[9][27] , \regfile[9][26] , \regfile[9][25] ,
         \regfile[9][24] , \regfile[9][23] , \regfile[9][22] ,
         \regfile[9][21] , \regfile[9][20] , \regfile[9][19] ,
         \regfile[9][18] , \regfile[9][17] , \regfile[9][16] ,
         \regfile[9][15] , \regfile[9][14] , \regfile[9][13] ,
         \regfile[9][12] , \regfile[9][11] , \regfile[9][10] , \regfile[9][9] ,
         \regfile[9][8] , \regfile[9][7] , \regfile[9][6] , \regfile[9][5] ,
         \regfile[9][4] , \regfile[9][3] , \regfile[9][2] , \regfile[9][1] ,
         \regfile[9][0] , \regfile[8][31] , \regfile[8][30] , \regfile[8][29] ,
         \regfile[8][28] , \regfile[8][27] , \regfile[8][26] ,
         \regfile[8][25] , \regfile[8][24] , \regfile[8][23] ,
         \regfile[8][22] , \regfile[8][21] , \regfile[8][20] ,
         \regfile[8][19] , \regfile[8][18] , \regfile[8][17] ,
         \regfile[8][16] , \regfile[8][15] , \regfile[8][14] ,
         \regfile[8][13] , \regfile[8][12] , \regfile[8][11] ,
         \regfile[8][10] , \regfile[8][9] , \regfile[8][8] , \regfile[8][7] ,
         \regfile[8][6] , \regfile[8][5] , \regfile[8][4] , \regfile[8][3] ,
         \regfile[8][2] , \regfile[8][1] , \regfile[8][0] , \regfile[7][31] ,
         \regfile[7][30] , \regfile[7][29] , \regfile[7][28] ,
         \regfile[7][27] , \regfile[7][26] , \regfile[7][25] ,
         \regfile[7][24] , \regfile[7][23] , \regfile[7][22] ,
         \regfile[7][21] , \regfile[7][20] , \regfile[7][19] ,
         \regfile[7][18] , \regfile[7][17] , \regfile[7][16] ,
         \regfile[7][15] , \regfile[7][14] , \regfile[7][13] ,
         \regfile[7][12] , \regfile[7][11] , \regfile[7][10] , \regfile[7][9] ,
         \regfile[7][8] , \regfile[7][7] , \regfile[7][6] , \regfile[7][5] ,
         \regfile[7][4] , \regfile[7][3] , \regfile[7][2] , \regfile[7][1] ,
         \regfile[7][0] , \regfile[6][31] , \regfile[6][30] , \regfile[6][29] ,
         \regfile[6][28] , \regfile[6][27] , \regfile[6][26] ,
         \regfile[6][25] , \regfile[6][24] , \regfile[6][23] ,
         \regfile[6][22] , \regfile[6][21] , \regfile[6][20] ,
         \regfile[6][19] , \regfile[6][18] , \regfile[6][17] ,
         \regfile[6][16] , \regfile[6][15] , \regfile[6][14] ,
         \regfile[6][13] , \regfile[6][12] , \regfile[6][11] ,
         \regfile[6][10] , \regfile[6][9] , \regfile[6][8] , \regfile[6][7] ,
         \regfile[6][6] , \regfile[6][5] , \regfile[6][4] , \regfile[6][3] ,
         \regfile[6][2] , \regfile[6][1] , \regfile[6][0] , \regfile[5][31] ,
         \regfile[5][30] , \regfile[5][29] , \regfile[5][28] ,
         \regfile[5][27] , \regfile[5][26] , \regfile[5][25] ,
         \regfile[5][24] , \regfile[5][23] , \regfile[5][22] ,
         \regfile[5][21] , \regfile[5][20] , \regfile[5][19] ,
         \regfile[5][18] , \regfile[5][17] , \regfile[5][16] ,
         \regfile[5][15] , \regfile[5][14] , \regfile[5][13] ,
         \regfile[5][12] , \regfile[5][11] , \regfile[5][10] , \regfile[5][9] ,
         \regfile[5][8] , \regfile[5][7] , \regfile[5][6] , \regfile[5][5] ,
         \regfile[5][4] , \regfile[5][3] , \regfile[5][2] , \regfile[5][1] ,
         \regfile[5][0] , \regfile[4][31] , \regfile[4][30] , \regfile[4][29] ,
         \regfile[4][28] , \regfile[4][27] , \regfile[4][26] ,
         \regfile[4][25] , \regfile[4][24] , \regfile[4][23] ,
         \regfile[4][22] , \regfile[4][21] , \regfile[4][20] ,
         \regfile[4][19] , \regfile[4][18] , \regfile[4][17] ,
         \regfile[4][16] , \regfile[4][15] , \regfile[4][14] ,
         \regfile[4][13] , \regfile[4][12] , \regfile[4][11] ,
         \regfile[4][10] , \regfile[4][9] , \regfile[4][8] , \regfile[4][7] ,
         \regfile[4][6] , \regfile[4][5] , \regfile[4][4] , \regfile[4][3] ,
         \regfile[4][2] , \regfile[4][1] , \regfile[4][0] , \regfile[3][31] ,
         \regfile[3][30] , \regfile[3][29] , \regfile[3][28] ,
         \regfile[3][27] , \regfile[3][26] , \regfile[3][25] ,
         \regfile[3][24] , \regfile[3][23] , \regfile[3][22] ,
         \regfile[3][21] , \regfile[3][20] , \regfile[3][19] ,
         \regfile[3][18] , \regfile[3][17] , \regfile[3][16] ,
         \regfile[3][15] , \regfile[3][14] , \regfile[3][13] ,
         \regfile[3][12] , \regfile[3][11] , \regfile[3][10] , \regfile[3][9] ,
         \regfile[3][8] , \regfile[3][7] , \regfile[3][6] , \regfile[3][5] ,
         \regfile[3][4] , \regfile[3][3] , \regfile[3][2] , \regfile[3][1] ,
         \regfile[3][0] , \regfile[2][31] , \regfile[2][30] , \regfile[2][29] ,
         \regfile[2][28] , \regfile[2][27] , \regfile[2][26] ,
         \regfile[2][25] , \regfile[2][24] , \regfile[2][23] ,
         \regfile[2][22] , \regfile[2][21] , \regfile[2][20] ,
         \regfile[2][19] , \regfile[2][18] , \regfile[2][17] ,
         \regfile[2][16] , \regfile[2][15] , \regfile[2][14] ,
         \regfile[2][13] , \regfile[2][12] , \regfile[2][11] ,
         \regfile[2][10] , \regfile[2][9] , \regfile[2][8] , \regfile[2][7] ,
         \regfile[2][6] , \regfile[2][5] , \regfile[2][4] , \regfile[2][3] ,
         \regfile[2][2] , \regfile[2][1] , \regfile[2][0] , \regfile[1][31] ,
         \regfile[1][30] , \regfile[1][29] , \regfile[1][28] ,
         \regfile[1][27] , \regfile[1][26] , \regfile[1][25] ,
         \regfile[1][24] , \regfile[1][23] , \regfile[1][22] ,
         \regfile[1][21] , \regfile[1][20] , \regfile[1][19] ,
         \regfile[1][18] , \regfile[1][17] , \regfile[1][16] ,
         \regfile[1][15] , \regfile[1][14] , \regfile[1][13] ,
         \regfile[1][12] , \regfile[1][11] , \regfile[1][10] , \regfile[1][9] ,
         \regfile[1][8] , \regfile[1][7] , \regfile[1][6] , \regfile[1][5] ,
         \regfile[1][4] , \regfile[1][3] , \regfile[1][2] , \regfile[1][1] ,
         \regfile[1][0] , \regfile[0][31] , \regfile[0][30] , \regfile[0][29] ,
         \regfile[0][28] , \regfile[0][27] , \regfile[0][26] ,
         \regfile[0][25] , \regfile[0][24] , \regfile[0][23] ,
         \regfile[0][22] , \regfile[0][21] , \regfile[0][20] ,
         \regfile[0][19] , \regfile[0][18] , \regfile[0][17] ,
         \regfile[0][16] , \regfile[0][15] , \regfile[0][14] ,
         \regfile[0][13] , \regfile[0][12] , \regfile[0][11] ,
         \regfile[0][10] , \regfile[0][9] , \regfile[0][8] , \regfile[0][7] ,
         \regfile[0][6] , \regfile[0][5] , \regfile[0][4] , \regfile[0][3] ,
         \regfile[0][2] , \regfile[0][1] , \regfile[0][0] , N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N254, N255, N256, N257, N258, N259, N260, N261,
         N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272,
         N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283,
         N284, N285, N286, N288, N289, N290, N291, N292, N293, N294, N295,
         N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306,
         N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317,
         N318, N319, N320, N321, N322, n10, n11, n12, n14, n15, n17, n18, n19,
         n21, n22, n24, n26, n29, n30, n32, n34, n36, n37, n39, n41, n44, n46,
         n48, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n66, n67,
         n68, n70, n72, n73, n75, n76, n77, n78, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n179, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172;
  wire   [3:0] opcode;
  wire   [31:0] tempA;
  wire   [31:0] tempB;
  assign N17 = instr[8];
  assign N18 = instr[9];
  assign N19 = instr[10];
  assign N20 = instr[11];
  assign N21 = instr[4];
  assign N22 = instr[5];
  assign N23 = instr[6];
  assign N24 = instr[7];

  DFFX1 \tempB_reg[31]  ( .D(N57), .CLK(clk), .Q(tempB[31]), .QN(n712) );
  DFFX1 \tempB_reg[30]  ( .D(N58), .CLK(clk), .Q(tempB[30]) );
  DFFX1 \tempB_reg[29]  ( .D(N59), .CLK(clk), .Q(tempB[29]) );
  DFFX1 \tempB_reg[28]  ( .D(N60), .CLK(clk), .Q(tempB[28]) );
  DFFX1 \tempB_reg[27]  ( .D(N61), .CLK(clk), .Q(tempB[27]) );
  DFFX1 \tempB_reg[26]  ( .D(N62), .CLK(clk), .Q(tempB[26]) );
  DFFX1 \tempB_reg[25]  ( .D(N63), .CLK(clk), .Q(tempB[25]) );
  DFFX1 \tempB_reg[24]  ( .D(N64), .CLK(clk), .Q(tempB[24]) );
  DFFX1 \tempB_reg[23]  ( .D(N65), .CLK(clk), .Q(tempB[23]) );
  DFFX1 \tempB_reg[22]  ( .D(N66), .CLK(clk), .Q(tempB[22]) );
  DFFX1 \tempB_reg[21]  ( .D(N67), .CLK(clk), .Q(tempB[21]) );
  DFFX1 \tempB_reg[20]  ( .D(N68), .CLK(clk), .Q(tempB[20]) );
  DFFX1 \tempB_reg[19]  ( .D(N69), .CLK(clk), .Q(tempB[19]) );
  DFFX1 \tempB_reg[18]  ( .D(N70), .CLK(clk), .Q(tempB[18]) );
  DFFX1 \tempB_reg[17]  ( .D(N71), .CLK(clk), .Q(tempB[17]) );
  DFFX1 \tempB_reg[16]  ( .D(N72), .CLK(clk), .Q(tempB[16]) );
  DFFX1 \tempB_reg[15]  ( .D(N73), .CLK(clk), .Q(tempB[15]) );
  DFFX1 \tempB_reg[14]  ( .D(N74), .CLK(clk), .Q(tempB[14]) );
  DFFX1 \tempB_reg[13]  ( .D(N75), .CLK(clk), .Q(tempB[13]) );
  DFFX1 \tempB_reg[12]  ( .D(N76), .CLK(clk), .Q(tempB[12]) );
  DFFX1 \tempB_reg[11]  ( .D(N77), .CLK(clk), .Q(tempB[11]) );
  DFFX1 \tempB_reg[10]  ( .D(N78), .CLK(clk), .Q(tempB[10]) );
  DFFX1 \tempB_reg[9]  ( .D(N79), .CLK(clk), .Q(tempB[9]) );
  DFFX1 \tempB_reg[8]  ( .D(N80), .CLK(clk), .Q(tempB[8]) );
  DFFX1 \tempB_reg[7]  ( .D(N81), .CLK(clk), .Q(tempB[7]) );
  DFFX1 \tempB_reg[6]  ( .D(N82), .CLK(clk), .Q(tempB[6]) );
  DFFX1 \tempB_reg[5]  ( .D(N83), .CLK(clk), .Q(tempB[5]) );
  DFFX1 \tempB_reg[4]  ( .D(N84), .CLK(clk), .Q(tempB[4]) );
  DFFX1 \tempB_reg[3]  ( .D(N85), .CLK(clk), .Q(tempB[3]) );
  DFFX1 \tempB_reg[2]  ( .D(N86), .CLK(clk), .Q(tempB[2]) );
  DFFX1 \tempB_reg[1]  ( .D(N87), .CLK(clk), .Q(tempB[1]) );
  DFFX1 \tempB_reg[0]  ( .D(N88), .CLK(clk), .Q(tempB[0]), .QN(n705) );
  DFFX1 \dest_reg[3]  ( .D(instr[3]), .CLK(clk), .Q(n704), .QN(n185) );
  DFFX1 \dest_reg[2]  ( .D(instr[2]), .CLK(clk), .Q(n708), .QN(n184) );
  DFFX1 \dest_reg[1]  ( .D(instr[1]), .CLK(clk), .Q(n709), .QN(n187) );
  DFFX1 \dest_reg[0]  ( .D(instr[0]), .CLK(clk), .Q(n703), .QN(n186) );
  DFFX1 \opcode_reg[3]  ( .D(instr[15]), .CLK(clk), .Q(opcode[3]) );
  DFFX1 \opcode_reg[2]  ( .D(instr[14]), .CLK(clk), .Q(n702), .QN(n700) );
  DFFX1 \opcode_reg[1]  ( .D(instr[13]), .CLK(clk), .Q(opcode[1]), .QN(n711)
         );
  DFFX1 \opcode_reg[0]  ( .D(instr[12]), .CLK(clk), .Q(n183), .QN(n706) );
  DFFX1 \tempA_reg[31]  ( .D(N25), .CLK(clk), .Q(tempA[31]), .QN(n707) );
  DFFX1 \tempA_reg[30]  ( .D(N26), .CLK(clk), .Q(tempA[30]) );
  DFFX1 \tempA_reg[29]  ( .D(N27), .CLK(clk), .Q(tempA[29]) );
  DFFX1 \tempA_reg[28]  ( .D(N28), .CLK(clk), .Q(tempA[28]) );
  DFFX1 \tempA_reg[27]  ( .D(N29), .CLK(clk), .Q(tempA[27]) );
  DFFX1 \tempA_reg[26]  ( .D(N30), .CLK(clk), .Q(tempA[26]) );
  DFFX1 \tempA_reg[25]  ( .D(N31), .CLK(clk), .Q(tempA[25]) );
  DFFX1 \tempA_reg[24]  ( .D(N32), .CLK(clk), .Q(tempA[24]) );
  DFFX1 \tempA_reg[23]  ( .D(N33), .CLK(clk), .Q(tempA[23]) );
  DFFX1 \tempA_reg[22]  ( .D(N34), .CLK(clk), .Q(tempA[22]) );
  DFFX1 \tempA_reg[21]  ( .D(N35), .CLK(clk), .Q(tempA[21]) );
  DFFX1 \tempA_reg[20]  ( .D(N36), .CLK(clk), .Q(tempA[20]) );
  DFFX1 \tempA_reg[19]  ( .D(N37), .CLK(clk), .Q(tempA[19]) );
  DFFX1 \tempA_reg[18]  ( .D(N38), .CLK(clk), .Q(tempA[18]) );
  DFFX1 \tempA_reg[17]  ( .D(N39), .CLK(clk), .Q(tempA[17]) );
  DFFX1 \tempA_reg[16]  ( .D(N40), .CLK(clk), .Q(tempA[16]) );
  DFFX1 \tempA_reg[15]  ( .D(N41), .CLK(clk), .Q(tempA[15]) );
  DFFX1 \tempA_reg[14]  ( .D(N42), .CLK(clk), .Q(tempA[14]) );
  DFFX1 \tempA_reg[13]  ( .D(N43), .CLK(clk), .Q(tempA[13]) );
  DFFX1 \tempA_reg[12]  ( .D(N44), .CLK(clk), .Q(tempA[12]) );
  DFFX1 \tempA_reg[11]  ( .D(N45), .CLK(clk), .Q(tempA[11]) );
  DFFX1 \tempA_reg[10]  ( .D(N46), .CLK(clk), .Q(tempA[10]) );
  DFFX1 \tempA_reg[9]  ( .D(N47), .CLK(clk), .Q(tempA[9]) );
  DFFX1 \tempA_reg[8]  ( .D(N48), .CLK(clk), .Q(tempA[8]) );
  DFFX1 \tempA_reg[7]  ( .D(N49), .CLK(clk), .Q(tempA[7]) );
  DFFX1 \tempA_reg[6]  ( .D(N50), .CLK(clk), .Q(tempA[6]) );
  DFFX1 \tempA_reg[5]  ( .D(N51), .CLK(clk), .Q(tempA[5]) );
  DFFX1 \tempA_reg[4]  ( .D(N52), .CLK(clk), .Q(tempA[4]) );
  DFFX1 \tempA_reg[3]  ( .D(N53), .CLK(clk), .Q(tempA[3]) );
  DFFX1 \tempA_reg[2]  ( .D(N54), .CLK(clk), .Q(tempA[2]) );
  DFFX1 \tempA_reg[1]  ( .D(N55), .CLK(clk), .Q(tempA[1]) );
  DFFX1 \tempA_reg[0]  ( .D(N56), .CLK(clk), .Q(tempA[0]), .QN(n710) );
  DFFX1 Overflow_reg ( .D(N322), .CLK(clk), .Q(Overflow) );
  DFFX1 \AluOut_reg[31]  ( .D(N321), .CLK(clk), .Q(AluOut[31]) );
  DFFX1 \AluOut_reg[30]  ( .D(N320), .CLK(clk), .Q(AluOut[30]) );
  DFFX1 \AluOut_reg[29]  ( .D(N319), .CLK(clk), .Q(AluOut[29]) );
  DFFX1 \AluOut_reg[28]  ( .D(N318), .CLK(clk), .Q(AluOut[28]) );
  DFFX1 \AluOut_reg[27]  ( .D(N317), .CLK(clk), .Q(AluOut[27]) );
  DFFX1 \AluOut_reg[26]  ( .D(N316), .CLK(clk), .Q(AluOut[26]) );
  DFFX1 \AluOut_reg[25]  ( .D(N315), .CLK(clk), .Q(AluOut[25]) );
  DFFX1 \AluOut_reg[24]  ( .D(N314), .CLK(clk), .Q(AluOut[24]) );
  DFFX1 \AluOut_reg[23]  ( .D(N313), .CLK(clk), .Q(AluOut[23]) );
  DFFX1 \AluOut_reg[22]  ( .D(N312), .CLK(clk), .Q(AluOut[22]) );
  DFFX1 \AluOut_reg[21]  ( .D(N311), .CLK(clk), .Q(AluOut[21]) );
  DFFX1 \AluOut_reg[20]  ( .D(N310), .CLK(clk), .Q(AluOut[20]) );
  DFFX1 \AluOut_reg[19]  ( .D(N309), .CLK(clk), .Q(AluOut[19]) );
  DFFX1 \AluOut_reg[18]  ( .D(N308), .CLK(clk), .Q(AluOut[18]) );
  DFFX1 \AluOut_reg[17]  ( .D(N307), .CLK(clk), .Q(AluOut[17]) );
  DFFX1 \AluOut_reg[16]  ( .D(N306), .CLK(clk), .Q(AluOut[16]) );
  DFFX1 \AluOut_reg[15]  ( .D(N305), .CLK(clk), .Q(AluOut[15]) );
  DFFX1 \AluOut_reg[14]  ( .D(N304), .CLK(clk), .Q(AluOut[14]) );
  DFFX1 \AluOut_reg[13]  ( .D(N303), .CLK(clk), .Q(AluOut[13]) );
  DFFX1 \AluOut_reg[12]  ( .D(N302), .CLK(clk), .Q(AluOut[12]) );
  DFFX1 \AluOut_reg[11]  ( .D(N301), .CLK(clk), .Q(AluOut[11]) );
  DFFX1 \AluOut_reg[10]  ( .D(N300), .CLK(clk), .Q(AluOut[10]) );
  DFFX1 \AluOut_reg[9]  ( .D(N299), .CLK(clk), .Q(AluOut[9]) );
  DFFX1 \AluOut_reg[8]  ( .D(N298), .CLK(clk), .Q(AluOut[8]) );
  DFFX1 \AluOut_reg[7]  ( .D(N297), .CLK(clk), .Q(AluOut[7]) );
  DFFX1 \AluOut_reg[6]  ( .D(N296), .CLK(clk), .Q(AluOut[6]) );
  DFFX1 \AluOut_reg[5]  ( .D(N295), .CLK(clk), .Q(AluOut[5]) );
  DFFX1 \AluOut_reg[4]  ( .D(N294), .CLK(clk), .Q(AluOut[4]) );
  DFFX1 \AluOut_reg[3]  ( .D(N293), .CLK(clk), .Q(AluOut[3]) );
  DFFX1 \AluOut_reg[2]  ( .D(N292), .CLK(clk), .Q(AluOut[2]) );
  DFFX1 \AluOut_reg[1]  ( .D(N291), .CLK(clk), .Q(AluOut[1]) );
  DFFX1 \AluOut_reg[0]  ( .D(N290), .CLK(clk), .Q(AluOut[0]) );
  DFFX1 Carryout_reg ( .D(N289), .CLK(clk), .Q(Carryout) );
  DFFX1 Zero_reg ( .D(n701), .CLK(clk), .Q(Zero) );
  DFFX1 \regfile_reg[15][31]  ( .D(n699), .CLK(clk), .Q(\regfile[15][31] ) );
  DFFX1 \regfile_reg[15][30]  ( .D(n698), .CLK(clk), .Q(\regfile[15][30] ) );
  DFFX1 \regfile_reg[15][29]  ( .D(n697), .CLK(clk), .Q(\regfile[15][29] ) );
  DFFX1 \regfile_reg[15][28]  ( .D(n696), .CLK(clk), .Q(\regfile[15][28] ) );
  DFFX1 \regfile_reg[15][27]  ( .D(n695), .CLK(clk), .Q(\regfile[15][27] ) );
  DFFX1 \regfile_reg[15][26]  ( .D(n694), .CLK(clk), .Q(\regfile[15][26] ) );
  DFFX1 \regfile_reg[15][25]  ( .D(n693), .CLK(clk), .Q(\regfile[15][25] ) );
  DFFX1 \regfile_reg[15][24]  ( .D(n692), .CLK(clk), .Q(\regfile[15][24] ) );
  DFFX1 \regfile_reg[15][23]  ( .D(n691), .CLK(clk), .Q(\regfile[15][23] ) );
  DFFX1 \regfile_reg[15][22]  ( .D(n690), .CLK(clk), .Q(\regfile[15][22] ) );
  DFFX1 \regfile_reg[15][21]  ( .D(n689), .CLK(clk), .Q(\regfile[15][21] ) );
  DFFX1 \regfile_reg[15][20]  ( .D(n688), .CLK(clk), .Q(\regfile[15][20] ) );
  DFFX1 \regfile_reg[15][19]  ( .D(n687), .CLK(clk), .Q(\regfile[15][19] ) );
  DFFX1 \regfile_reg[15][18]  ( .D(n686), .CLK(clk), .Q(\regfile[15][18] ) );
  DFFX1 \regfile_reg[15][17]  ( .D(n685), .CLK(clk), .Q(\regfile[15][17] ) );
  DFFX1 \regfile_reg[15][16]  ( .D(n684), .CLK(clk), .Q(\regfile[15][16] ) );
  DFFX1 \regfile_reg[15][15]  ( .D(n683), .CLK(clk), .Q(\regfile[15][15] ) );
  DFFX1 \regfile_reg[15][14]  ( .D(n682), .CLK(clk), .Q(\regfile[15][14] ) );
  DFFX1 \regfile_reg[15][13]  ( .D(n681), .CLK(clk), .Q(\regfile[15][13] ) );
  DFFX1 \regfile_reg[15][12]  ( .D(n680), .CLK(clk), .Q(\regfile[15][12] ) );
  DFFX1 \regfile_reg[15][11]  ( .D(n679), .CLK(clk), .Q(\regfile[15][11] ) );
  DFFX1 \regfile_reg[15][10]  ( .D(n678), .CLK(clk), .Q(\regfile[15][10] ) );
  DFFX1 \regfile_reg[15][9]  ( .D(n677), .CLK(clk), .Q(\regfile[15][9] ) );
  DFFX1 \regfile_reg[15][8]  ( .D(n676), .CLK(clk), .Q(\regfile[15][8] ) );
  DFFX1 \regfile_reg[15][7]  ( .D(n675), .CLK(clk), .Q(\regfile[15][7] ) );
  DFFX1 \regfile_reg[15][6]  ( .D(n674), .CLK(clk), .Q(\regfile[15][6] ) );
  DFFX1 \regfile_reg[15][5]  ( .D(n673), .CLK(clk), .Q(\regfile[15][5] ) );
  DFFX1 \regfile_reg[15][4]  ( .D(n672), .CLK(clk), .Q(\regfile[15][4] ) );
  DFFX1 \regfile_reg[15][3]  ( .D(n671), .CLK(clk), .Q(\regfile[15][3] ) );
  DFFX1 \regfile_reg[15][2]  ( .D(n670), .CLK(clk), .Q(\regfile[15][2] ) );
  DFFX1 \regfile_reg[15][1]  ( .D(n669), .CLK(clk), .Q(\regfile[15][1] ) );
  DFFX1 \regfile_reg[15][0]  ( .D(n668), .CLK(clk), .Q(\regfile[15][0] ) );
  DFFX1 \regfile_reg[14][31]  ( .D(n667), .CLK(clk), .Q(\regfile[14][31] ) );
  DFFX1 \regfile_reg[14][30]  ( .D(n666), .CLK(clk), .Q(\regfile[14][30] ) );
  DFFX1 \regfile_reg[14][29]  ( .D(n665), .CLK(clk), .Q(\regfile[14][29] ) );
  DFFX1 \regfile_reg[14][28]  ( .D(n664), .CLK(clk), .Q(\regfile[14][28] ) );
  DFFX1 \regfile_reg[14][27]  ( .D(n663), .CLK(clk), .Q(\regfile[14][27] ) );
  DFFX1 \regfile_reg[14][26]  ( .D(n662), .CLK(clk), .Q(\regfile[14][26] ) );
  DFFX1 \regfile_reg[14][25]  ( .D(n661), .CLK(clk), .Q(\regfile[14][25] ) );
  DFFX1 \regfile_reg[14][24]  ( .D(n660), .CLK(clk), .Q(\regfile[14][24] ) );
  DFFX1 \regfile_reg[14][23]  ( .D(n659), .CLK(clk), .Q(\regfile[14][23] ) );
  DFFX1 \regfile_reg[14][22]  ( .D(n658), .CLK(clk), .Q(\regfile[14][22] ) );
  DFFX1 \regfile_reg[14][21]  ( .D(n657), .CLK(clk), .Q(\regfile[14][21] ) );
  DFFX1 \regfile_reg[14][20]  ( .D(n656), .CLK(clk), .Q(\regfile[14][20] ) );
  DFFX1 \regfile_reg[14][19]  ( .D(n655), .CLK(clk), .Q(\regfile[14][19] ) );
  DFFX1 \regfile_reg[14][18]  ( .D(n654), .CLK(clk), .Q(\regfile[14][18] ) );
  DFFX1 \regfile_reg[14][17]  ( .D(n653), .CLK(clk), .Q(\regfile[14][17] ) );
  DFFX1 \regfile_reg[14][16]  ( .D(n652), .CLK(clk), .Q(\regfile[14][16] ) );
  DFFX1 \regfile_reg[14][15]  ( .D(n651), .CLK(clk), .Q(\regfile[14][15] ) );
  DFFX1 \regfile_reg[14][14]  ( .D(n650), .CLK(clk), .Q(\regfile[14][14] ) );
  DFFX1 \regfile_reg[14][13]  ( .D(n649), .CLK(clk), .Q(\regfile[14][13] ) );
  DFFX1 \regfile_reg[14][12]  ( .D(n648), .CLK(clk), .Q(\regfile[14][12] ) );
  DFFX1 \regfile_reg[14][11]  ( .D(n647), .CLK(clk), .Q(\regfile[14][11] ) );
  DFFX1 \regfile_reg[14][10]  ( .D(n646), .CLK(clk), .Q(\regfile[14][10] ) );
  DFFX1 \regfile_reg[14][9]  ( .D(n645), .CLK(clk), .Q(\regfile[14][9] ) );
  DFFX1 \regfile_reg[14][8]  ( .D(n644), .CLK(clk), .Q(\regfile[14][8] ) );
  DFFX1 \regfile_reg[14][7]  ( .D(n643), .CLK(clk), .Q(\regfile[14][7] ) );
  DFFX1 \regfile_reg[14][6]  ( .D(n642), .CLK(clk), .Q(\regfile[14][6] ) );
  DFFX1 \regfile_reg[14][5]  ( .D(n641), .CLK(clk), .Q(\regfile[14][5] ) );
  DFFX1 \regfile_reg[14][4]  ( .D(n640), .CLK(clk), .Q(\regfile[14][4] ) );
  DFFX1 \regfile_reg[14][3]  ( .D(n639), .CLK(clk), .Q(\regfile[14][3] ) );
  DFFX1 \regfile_reg[14][2]  ( .D(n638), .CLK(clk), .Q(\regfile[14][2] ) );
  DFFX1 \regfile_reg[14][1]  ( .D(n637), .CLK(clk), .Q(\regfile[14][1] ) );
  DFFX1 \regfile_reg[14][0]  ( .D(n636), .CLK(clk), .Q(\regfile[14][0] ) );
  DFFX1 \regfile_reg[13][31]  ( .D(n635), .CLK(clk), .Q(\regfile[13][31] ) );
  DFFX1 \regfile_reg[13][30]  ( .D(n634), .CLK(clk), .Q(\regfile[13][30] ) );
  DFFX1 \regfile_reg[13][29]  ( .D(n633), .CLK(clk), .Q(\regfile[13][29] ) );
  DFFX1 \regfile_reg[13][28]  ( .D(n632), .CLK(clk), .Q(\regfile[13][28] ) );
  DFFX1 \regfile_reg[13][27]  ( .D(n631), .CLK(clk), .Q(\regfile[13][27] ) );
  DFFX1 \regfile_reg[13][26]  ( .D(n630), .CLK(clk), .Q(\regfile[13][26] ) );
  DFFX1 \regfile_reg[13][25]  ( .D(n629), .CLK(clk), .Q(\regfile[13][25] ) );
  DFFX1 \regfile_reg[13][24]  ( .D(n628), .CLK(clk), .Q(\regfile[13][24] ) );
  DFFX1 \regfile_reg[13][23]  ( .D(n627), .CLK(clk), .Q(\regfile[13][23] ) );
  DFFX1 \regfile_reg[13][22]  ( .D(n626), .CLK(clk), .Q(\regfile[13][22] ) );
  DFFX1 \regfile_reg[13][21]  ( .D(n625), .CLK(clk), .Q(\regfile[13][21] ) );
  DFFX1 \regfile_reg[13][20]  ( .D(n624), .CLK(clk), .Q(\regfile[13][20] ) );
  DFFX1 \regfile_reg[13][19]  ( .D(n623), .CLK(clk), .Q(\regfile[13][19] ) );
  DFFX1 \regfile_reg[13][18]  ( .D(n622), .CLK(clk), .Q(\regfile[13][18] ) );
  DFFX1 \regfile_reg[13][17]  ( .D(n621), .CLK(clk), .Q(\regfile[13][17] ) );
  DFFX1 \regfile_reg[13][16]  ( .D(n620), .CLK(clk), .Q(\regfile[13][16] ) );
  DFFX1 \regfile_reg[13][15]  ( .D(n619), .CLK(clk), .Q(\regfile[13][15] ) );
  DFFX1 \regfile_reg[13][14]  ( .D(n618), .CLK(clk), .Q(\regfile[13][14] ) );
  DFFX1 \regfile_reg[13][13]  ( .D(n617), .CLK(clk), .Q(\regfile[13][13] ) );
  DFFX1 \regfile_reg[13][12]  ( .D(n616), .CLK(clk), .Q(\regfile[13][12] ) );
  DFFX1 \regfile_reg[13][11]  ( .D(n615), .CLK(clk), .Q(\regfile[13][11] ) );
  DFFX1 \regfile_reg[13][10]  ( .D(n614), .CLK(clk), .Q(\regfile[13][10] ) );
  DFFX1 \regfile_reg[13][9]  ( .D(n613), .CLK(clk), .Q(\regfile[13][9] ) );
  DFFX1 \regfile_reg[13][8]  ( .D(n612), .CLK(clk), .Q(\regfile[13][8] ) );
  DFFX1 \regfile_reg[13][7]  ( .D(n611), .CLK(clk), .Q(\regfile[13][7] ) );
  DFFX1 \regfile_reg[13][6]  ( .D(n610), .CLK(clk), .Q(\regfile[13][6] ) );
  DFFX1 \regfile_reg[13][5]  ( .D(n609), .CLK(clk), .Q(\regfile[13][5] ) );
  DFFX1 \regfile_reg[13][4]  ( .D(n608), .CLK(clk), .Q(\regfile[13][4] ) );
  DFFX1 \regfile_reg[13][3]  ( .D(n607), .CLK(clk), .Q(\regfile[13][3] ) );
  DFFX1 \regfile_reg[13][2]  ( .D(n606), .CLK(clk), .Q(\regfile[13][2] ) );
  DFFX1 \regfile_reg[13][1]  ( .D(n605), .CLK(clk), .Q(\regfile[13][1] ) );
  DFFX1 \regfile_reg[13][0]  ( .D(n604), .CLK(clk), .Q(\regfile[13][0] ) );
  DFFX1 \regfile_reg[12][31]  ( .D(n603), .CLK(clk), .Q(\regfile[12][31] ) );
  DFFX1 \regfile_reg[12][30]  ( .D(n602), .CLK(clk), .Q(\regfile[12][30] ) );
  DFFX1 \regfile_reg[12][29]  ( .D(n601), .CLK(clk), .Q(\regfile[12][29] ) );
  DFFX1 \regfile_reg[12][28]  ( .D(n600), .CLK(clk), .Q(\regfile[12][28] ) );
  DFFX1 \regfile_reg[12][27]  ( .D(n599), .CLK(clk), .Q(\regfile[12][27] ) );
  DFFX1 \regfile_reg[12][26]  ( .D(n598), .CLK(clk), .Q(\regfile[12][26] ) );
  DFFX1 \regfile_reg[12][25]  ( .D(n597), .CLK(clk), .Q(\regfile[12][25] ) );
  DFFX1 \regfile_reg[12][24]  ( .D(n596), .CLK(clk), .Q(\regfile[12][24] ) );
  DFFX1 \regfile_reg[12][23]  ( .D(n595), .CLK(clk), .Q(\regfile[12][23] ) );
  DFFX1 \regfile_reg[12][22]  ( .D(n594), .CLK(clk), .Q(\regfile[12][22] ) );
  DFFX1 \regfile_reg[12][21]  ( .D(n593), .CLK(clk), .Q(\regfile[12][21] ) );
  DFFX1 \regfile_reg[12][20]  ( .D(n592), .CLK(clk), .Q(\regfile[12][20] ) );
  DFFX1 \regfile_reg[12][19]  ( .D(n591), .CLK(clk), .Q(\regfile[12][19] ) );
  DFFX1 \regfile_reg[12][18]  ( .D(n590), .CLK(clk), .Q(\regfile[12][18] ) );
  DFFX1 \regfile_reg[12][17]  ( .D(n589), .CLK(clk), .Q(\regfile[12][17] ) );
  DFFX1 \regfile_reg[12][16]  ( .D(n588), .CLK(clk), .Q(\regfile[12][16] ) );
  DFFX1 \regfile_reg[12][15]  ( .D(n587), .CLK(clk), .Q(\regfile[12][15] ) );
  DFFX1 \regfile_reg[12][14]  ( .D(n586), .CLK(clk), .Q(\regfile[12][14] ) );
  DFFX1 \regfile_reg[12][13]  ( .D(n585), .CLK(clk), .Q(\regfile[12][13] ) );
  DFFX1 \regfile_reg[12][12]  ( .D(n584), .CLK(clk), .Q(\regfile[12][12] ) );
  DFFX1 \regfile_reg[12][11]  ( .D(n583), .CLK(clk), .Q(\regfile[12][11] ) );
  DFFX1 \regfile_reg[12][10]  ( .D(n582), .CLK(clk), .Q(\regfile[12][10] ) );
  DFFX1 \regfile_reg[12][9]  ( .D(n581), .CLK(clk), .Q(\regfile[12][9] ) );
  DFFX1 \regfile_reg[12][8]  ( .D(n580), .CLK(clk), .Q(\regfile[12][8] ) );
  DFFX1 \regfile_reg[12][7]  ( .D(n579), .CLK(clk), .Q(\regfile[12][7] ) );
  DFFX1 \regfile_reg[12][6]  ( .D(n578), .CLK(clk), .Q(\regfile[12][6] ) );
  DFFX1 \regfile_reg[12][5]  ( .D(n577), .CLK(clk), .Q(\regfile[12][5] ) );
  DFFX1 \regfile_reg[12][4]  ( .D(n576), .CLK(clk), .Q(\regfile[12][4] ) );
  DFFX1 \regfile_reg[12][3]  ( .D(n575), .CLK(clk), .Q(\regfile[12][3] ) );
  DFFX1 \regfile_reg[12][2]  ( .D(n574), .CLK(clk), .Q(\regfile[12][2] ) );
  DFFX1 \regfile_reg[12][1]  ( .D(n573), .CLK(clk), .Q(\regfile[12][1] ) );
  DFFX1 \regfile_reg[12][0]  ( .D(n572), .CLK(clk), .Q(\regfile[12][0] ) );
  DFFX1 \regfile_reg[11][31]  ( .D(n571), .CLK(clk), .Q(\regfile[11][31] ) );
  DFFX1 \regfile_reg[11][30]  ( .D(n570), .CLK(clk), .Q(\regfile[11][30] ) );
  DFFX1 \regfile_reg[11][29]  ( .D(n569), .CLK(clk), .Q(\regfile[11][29] ) );
  DFFX1 \regfile_reg[11][28]  ( .D(n568), .CLK(clk), .Q(\regfile[11][28] ) );
  DFFX1 \regfile_reg[11][27]  ( .D(n567), .CLK(clk), .Q(\regfile[11][27] ) );
  DFFX1 \regfile_reg[11][26]  ( .D(n566), .CLK(clk), .Q(\regfile[11][26] ) );
  DFFX1 \regfile_reg[11][25]  ( .D(n565), .CLK(clk), .Q(\regfile[11][25] ) );
  DFFX1 \regfile_reg[11][24]  ( .D(n564), .CLK(clk), .Q(\regfile[11][24] ) );
  DFFX1 \regfile_reg[11][23]  ( .D(n563), .CLK(clk), .Q(\regfile[11][23] ) );
  DFFX1 \regfile_reg[11][22]  ( .D(n562), .CLK(clk), .Q(\regfile[11][22] ) );
  DFFX1 \regfile_reg[11][21]  ( .D(n561), .CLK(clk), .Q(\regfile[11][21] ) );
  DFFX1 \regfile_reg[11][20]  ( .D(n560), .CLK(clk), .Q(\regfile[11][20] ) );
  DFFX1 \regfile_reg[11][19]  ( .D(n559), .CLK(clk), .Q(\regfile[11][19] ) );
  DFFX1 \regfile_reg[11][18]  ( .D(n558), .CLK(clk), .Q(\regfile[11][18] ) );
  DFFX1 \regfile_reg[11][17]  ( .D(n557), .CLK(clk), .Q(\regfile[11][17] ) );
  DFFX1 \regfile_reg[11][16]  ( .D(n556), .CLK(clk), .Q(\regfile[11][16] ) );
  DFFX1 \regfile_reg[11][15]  ( .D(n555), .CLK(clk), .Q(\regfile[11][15] ) );
  DFFX1 \regfile_reg[11][14]  ( .D(n554), .CLK(clk), .Q(\regfile[11][14] ) );
  DFFX1 \regfile_reg[11][13]  ( .D(n553), .CLK(clk), .Q(\regfile[11][13] ) );
  DFFX1 \regfile_reg[11][12]  ( .D(n552), .CLK(clk), .Q(\regfile[11][12] ) );
  DFFX1 \regfile_reg[11][11]  ( .D(n551), .CLK(clk), .Q(\regfile[11][11] ) );
  DFFX1 \regfile_reg[11][10]  ( .D(n550), .CLK(clk), .Q(\regfile[11][10] ) );
  DFFX1 \regfile_reg[11][9]  ( .D(n549), .CLK(clk), .Q(\regfile[11][9] ) );
  DFFX1 \regfile_reg[11][8]  ( .D(n548), .CLK(clk), .Q(\regfile[11][8] ) );
  DFFX1 \regfile_reg[11][7]  ( .D(n547), .CLK(clk), .Q(\regfile[11][7] ) );
  DFFX1 \regfile_reg[11][6]  ( .D(n546), .CLK(clk), .Q(\regfile[11][6] ) );
  DFFX1 \regfile_reg[11][5]  ( .D(n545), .CLK(clk), .Q(\regfile[11][5] ) );
  DFFX1 \regfile_reg[11][4]  ( .D(n544), .CLK(clk), .Q(\regfile[11][4] ) );
  DFFX1 \regfile_reg[11][3]  ( .D(n543), .CLK(clk), .Q(\regfile[11][3] ) );
  DFFX1 \regfile_reg[11][2]  ( .D(n542), .CLK(clk), .Q(\regfile[11][2] ) );
  DFFX1 \regfile_reg[11][1]  ( .D(n541), .CLK(clk), .Q(\regfile[11][1] ) );
  DFFX1 \regfile_reg[11][0]  ( .D(n540), .CLK(clk), .Q(\regfile[11][0] ) );
  DFFX1 \regfile_reg[10][31]  ( .D(n539), .CLK(clk), .Q(\regfile[10][31] ) );
  DFFX1 \regfile_reg[10][30]  ( .D(n538), .CLK(clk), .Q(\regfile[10][30] ) );
  DFFX1 \regfile_reg[10][29]  ( .D(n537), .CLK(clk), .Q(\regfile[10][29] ) );
  DFFX1 \regfile_reg[10][28]  ( .D(n536), .CLK(clk), .Q(\regfile[10][28] ) );
  DFFX1 \regfile_reg[10][27]  ( .D(n535), .CLK(clk), .Q(\regfile[10][27] ) );
  DFFX1 \regfile_reg[10][26]  ( .D(n534), .CLK(clk), .Q(\regfile[10][26] ) );
  DFFX1 \regfile_reg[10][25]  ( .D(n533), .CLK(clk), .Q(\regfile[10][25] ) );
  DFFX1 \regfile_reg[10][24]  ( .D(n532), .CLK(clk), .Q(\regfile[10][24] ) );
  DFFX1 \regfile_reg[10][23]  ( .D(n531), .CLK(clk), .Q(\regfile[10][23] ) );
  DFFX1 \regfile_reg[10][22]  ( .D(n530), .CLK(clk), .Q(\regfile[10][22] ) );
  DFFX1 \regfile_reg[10][21]  ( .D(n529), .CLK(clk), .Q(\regfile[10][21] ) );
  DFFX1 \regfile_reg[10][20]  ( .D(n528), .CLK(clk), .Q(\regfile[10][20] ) );
  DFFX1 \regfile_reg[10][19]  ( .D(n527), .CLK(clk), .Q(\regfile[10][19] ) );
  DFFX1 \regfile_reg[10][18]  ( .D(n526), .CLK(clk), .Q(\regfile[10][18] ) );
  DFFX1 \regfile_reg[10][17]  ( .D(n525), .CLK(clk), .Q(\regfile[10][17] ) );
  DFFX1 \regfile_reg[10][16]  ( .D(n524), .CLK(clk), .Q(\regfile[10][16] ) );
  DFFX1 \regfile_reg[10][15]  ( .D(n523), .CLK(clk), .Q(\regfile[10][15] ) );
  DFFX1 \regfile_reg[10][14]  ( .D(n522), .CLK(clk), .Q(\regfile[10][14] ) );
  DFFX1 \regfile_reg[10][13]  ( .D(n521), .CLK(clk), .Q(\regfile[10][13] ) );
  DFFX1 \regfile_reg[10][12]  ( .D(n520), .CLK(clk), .Q(\regfile[10][12] ) );
  DFFX1 \regfile_reg[10][11]  ( .D(n519), .CLK(clk), .Q(\regfile[10][11] ) );
  DFFX1 \regfile_reg[10][10]  ( .D(n518), .CLK(clk), .Q(\regfile[10][10] ) );
  DFFX1 \regfile_reg[10][9]  ( .D(n517), .CLK(clk), .Q(\regfile[10][9] ) );
  DFFX1 \regfile_reg[10][8]  ( .D(n516), .CLK(clk), .Q(\regfile[10][8] ) );
  DFFX1 \regfile_reg[10][7]  ( .D(n515), .CLK(clk), .Q(\regfile[10][7] ) );
  DFFX1 \regfile_reg[10][6]  ( .D(n514), .CLK(clk), .Q(\regfile[10][6] ) );
  DFFX1 \regfile_reg[10][5]  ( .D(n513), .CLK(clk), .Q(\regfile[10][5] ) );
  DFFX1 \regfile_reg[10][4]  ( .D(n512), .CLK(clk), .Q(\regfile[10][4] ) );
  DFFX1 \regfile_reg[10][3]  ( .D(n511), .CLK(clk), .Q(\regfile[10][3] ) );
  DFFX1 \regfile_reg[10][2]  ( .D(n510), .CLK(clk), .Q(\regfile[10][2] ) );
  DFFX1 \regfile_reg[10][1]  ( .D(n509), .CLK(clk), .Q(\regfile[10][1] ) );
  DFFX1 \regfile_reg[10][0]  ( .D(n508), .CLK(clk), .Q(\regfile[10][0] ) );
  DFFX1 \regfile_reg[9][31]  ( .D(n507), .CLK(clk), .Q(\regfile[9][31] ) );
  DFFX1 \regfile_reg[9][30]  ( .D(n506), .CLK(clk), .Q(\regfile[9][30] ) );
  DFFX1 \regfile_reg[9][29]  ( .D(n505), .CLK(clk), .Q(\regfile[9][29] ) );
  DFFX1 \regfile_reg[9][28]  ( .D(n504), .CLK(clk), .Q(\regfile[9][28] ) );
  DFFX1 \regfile_reg[9][27]  ( .D(n503), .CLK(clk), .Q(\regfile[9][27] ) );
  DFFX1 \regfile_reg[9][26]  ( .D(n502), .CLK(clk), .Q(\regfile[9][26] ) );
  DFFX1 \regfile_reg[9][25]  ( .D(n501), .CLK(clk), .Q(\regfile[9][25] ) );
  DFFX1 \regfile_reg[9][24]  ( .D(n500), .CLK(clk), .Q(\regfile[9][24] ) );
  DFFX1 \regfile_reg[9][23]  ( .D(n499), .CLK(clk), .Q(\regfile[9][23] ) );
  DFFX1 \regfile_reg[9][22]  ( .D(n498), .CLK(clk), .Q(\regfile[9][22] ) );
  DFFX1 \regfile_reg[9][21]  ( .D(n497), .CLK(clk), .Q(\regfile[9][21] ) );
  DFFX1 \regfile_reg[9][20]  ( .D(n496), .CLK(clk), .Q(\regfile[9][20] ) );
  DFFX1 \regfile_reg[9][19]  ( .D(n495), .CLK(clk), .Q(\regfile[9][19] ) );
  DFFX1 \regfile_reg[9][18]  ( .D(n494), .CLK(clk), .Q(\regfile[9][18] ) );
  DFFX1 \regfile_reg[9][17]  ( .D(n493), .CLK(clk), .Q(\regfile[9][17] ) );
  DFFX1 \regfile_reg[9][16]  ( .D(n492), .CLK(clk), .Q(\regfile[9][16] ) );
  DFFX1 \regfile_reg[9][15]  ( .D(n491), .CLK(clk), .Q(\regfile[9][15] ) );
  DFFX1 \regfile_reg[9][14]  ( .D(n490), .CLK(clk), .Q(\regfile[9][14] ) );
  DFFX1 \regfile_reg[9][13]  ( .D(n489), .CLK(clk), .Q(\regfile[9][13] ) );
  DFFX1 \regfile_reg[9][12]  ( .D(n488), .CLK(clk), .Q(\regfile[9][12] ) );
  DFFX1 \regfile_reg[9][11]  ( .D(n487), .CLK(clk), .Q(\regfile[9][11] ) );
  DFFX1 \regfile_reg[9][10]  ( .D(n486), .CLK(clk), .Q(\regfile[9][10] ) );
  DFFX1 \regfile_reg[9][9]  ( .D(n485), .CLK(clk), .Q(\regfile[9][9] ) );
  DFFX1 \regfile_reg[9][8]  ( .D(n484), .CLK(clk), .Q(\regfile[9][8] ) );
  DFFX1 \regfile_reg[9][7]  ( .D(n483), .CLK(clk), .Q(\regfile[9][7] ) );
  DFFX1 \regfile_reg[9][6]  ( .D(n482), .CLK(clk), .Q(\regfile[9][6] ) );
  DFFX1 \regfile_reg[9][5]  ( .D(n481), .CLK(clk), .Q(\regfile[9][5] ) );
  DFFX1 \regfile_reg[9][4]  ( .D(n480), .CLK(clk), .Q(\regfile[9][4] ) );
  DFFX1 \regfile_reg[9][3]  ( .D(n479), .CLK(clk), .Q(\regfile[9][3] ) );
  DFFX1 \regfile_reg[9][2]  ( .D(n478), .CLK(clk), .Q(\regfile[9][2] ) );
  DFFX1 \regfile_reg[9][1]  ( .D(n477), .CLK(clk), .Q(\regfile[9][1] ) );
  DFFX1 \regfile_reg[9][0]  ( .D(n476), .CLK(clk), .Q(\regfile[9][0] ) );
  DFFX1 \regfile_reg[8][31]  ( .D(n475), .CLK(clk), .Q(\regfile[8][31] ) );
  DFFX1 \regfile_reg[8][30]  ( .D(n474), .CLK(clk), .Q(\regfile[8][30] ) );
  DFFX1 \regfile_reg[8][29]  ( .D(n473), .CLK(clk), .Q(\regfile[8][29] ) );
  DFFX1 \regfile_reg[8][28]  ( .D(n472), .CLK(clk), .Q(\regfile[8][28] ) );
  DFFX1 \regfile_reg[8][27]  ( .D(n471), .CLK(clk), .Q(\regfile[8][27] ) );
  DFFX1 \regfile_reg[8][26]  ( .D(n470), .CLK(clk), .Q(\regfile[8][26] ) );
  DFFX1 \regfile_reg[8][25]  ( .D(n469), .CLK(clk), .Q(\regfile[8][25] ) );
  DFFX1 \regfile_reg[8][24]  ( .D(n468), .CLK(clk), .Q(\regfile[8][24] ) );
  DFFX1 \regfile_reg[8][23]  ( .D(n467), .CLK(clk), .Q(\regfile[8][23] ) );
  DFFX1 \regfile_reg[8][22]  ( .D(n466), .CLK(clk), .Q(\regfile[8][22] ) );
  DFFX1 \regfile_reg[8][21]  ( .D(n465), .CLK(clk), .Q(\regfile[8][21] ) );
  DFFX1 \regfile_reg[8][20]  ( .D(n464), .CLK(clk), .Q(\regfile[8][20] ) );
  DFFX1 \regfile_reg[8][19]  ( .D(n463), .CLK(clk), .Q(\regfile[8][19] ) );
  DFFX1 \regfile_reg[8][18]  ( .D(n462), .CLK(clk), .Q(\regfile[8][18] ) );
  DFFX1 \regfile_reg[8][17]  ( .D(n461), .CLK(clk), .Q(\regfile[8][17] ) );
  DFFX1 \regfile_reg[8][16]  ( .D(n460), .CLK(clk), .Q(\regfile[8][16] ) );
  DFFX1 \regfile_reg[8][15]  ( .D(n459), .CLK(clk), .Q(\regfile[8][15] ) );
  DFFX1 \regfile_reg[8][14]  ( .D(n458), .CLK(clk), .Q(\regfile[8][14] ) );
  DFFX1 \regfile_reg[8][13]  ( .D(n457), .CLK(clk), .Q(\regfile[8][13] ) );
  DFFX1 \regfile_reg[8][12]  ( .D(n456), .CLK(clk), .Q(\regfile[8][12] ) );
  DFFX1 \regfile_reg[8][11]  ( .D(n455), .CLK(clk), .Q(\regfile[8][11] ) );
  DFFX1 \regfile_reg[8][10]  ( .D(n454), .CLK(clk), .Q(\regfile[8][10] ) );
  DFFX1 \regfile_reg[8][9]  ( .D(n453), .CLK(clk), .Q(\regfile[8][9] ) );
  DFFX1 \regfile_reg[8][8]  ( .D(n452), .CLK(clk), .Q(\regfile[8][8] ) );
  DFFX1 \regfile_reg[8][7]  ( .D(n451), .CLK(clk), .Q(\regfile[8][7] ) );
  DFFX1 \regfile_reg[8][6]  ( .D(n450), .CLK(clk), .Q(\regfile[8][6] ) );
  DFFX1 \regfile_reg[8][5]  ( .D(n449), .CLK(clk), .Q(\regfile[8][5] ) );
  DFFX1 \regfile_reg[8][4]  ( .D(n448), .CLK(clk), .Q(\regfile[8][4] ) );
  DFFX1 \regfile_reg[8][3]  ( .D(n447), .CLK(clk), .Q(\regfile[8][3] ) );
  DFFX1 \regfile_reg[8][2]  ( .D(n446), .CLK(clk), .Q(\regfile[8][2] ) );
  DFFX1 \regfile_reg[8][1]  ( .D(n445), .CLK(clk), .Q(\regfile[8][1] ) );
  DFFX1 \regfile_reg[8][0]  ( .D(n444), .CLK(clk), .Q(\regfile[8][0] ) );
  DFFX1 \regfile_reg[7][31]  ( .D(n443), .CLK(clk), .Q(\regfile[7][31] ) );
  DFFX1 \regfile_reg[7][30]  ( .D(n442), .CLK(clk), .Q(\regfile[7][30] ) );
  DFFX1 \regfile_reg[7][29]  ( .D(n441), .CLK(clk), .Q(\regfile[7][29] ) );
  DFFX1 \regfile_reg[7][28]  ( .D(n440), .CLK(clk), .Q(\regfile[7][28] ) );
  DFFX1 \regfile_reg[7][27]  ( .D(n439), .CLK(clk), .Q(\regfile[7][27] ) );
  DFFX1 \regfile_reg[7][26]  ( .D(n438), .CLK(clk), .Q(\regfile[7][26] ) );
  DFFX1 \regfile_reg[7][25]  ( .D(n437), .CLK(clk), .Q(\regfile[7][25] ) );
  DFFX1 \regfile_reg[7][24]  ( .D(n436), .CLK(clk), .Q(\regfile[7][24] ) );
  DFFX1 \regfile_reg[7][23]  ( .D(n435), .CLK(clk), .Q(\regfile[7][23] ) );
  DFFX1 \regfile_reg[7][22]  ( .D(n434), .CLK(clk), .Q(\regfile[7][22] ) );
  DFFX1 \regfile_reg[7][21]  ( .D(n433), .CLK(clk), .Q(\regfile[7][21] ) );
  DFFX1 \regfile_reg[7][20]  ( .D(n432), .CLK(clk), .Q(\regfile[7][20] ) );
  DFFX1 \regfile_reg[7][19]  ( .D(n431), .CLK(clk), .Q(\regfile[7][19] ) );
  DFFX1 \regfile_reg[7][18]  ( .D(n430), .CLK(clk), .Q(\regfile[7][18] ) );
  DFFX1 \regfile_reg[7][17]  ( .D(n429), .CLK(clk), .Q(\regfile[7][17] ) );
  DFFX1 \regfile_reg[7][16]  ( .D(n428), .CLK(clk), .Q(\regfile[7][16] ) );
  DFFX1 \regfile_reg[7][15]  ( .D(n427), .CLK(clk), .Q(\regfile[7][15] ) );
  DFFX1 \regfile_reg[7][14]  ( .D(n426), .CLK(clk), .Q(\regfile[7][14] ) );
  DFFX1 \regfile_reg[7][13]  ( .D(n425), .CLK(clk), .Q(\regfile[7][13] ) );
  DFFX1 \regfile_reg[7][12]  ( .D(n424), .CLK(clk), .Q(\regfile[7][12] ) );
  DFFX1 \regfile_reg[7][11]  ( .D(n423), .CLK(clk), .Q(\regfile[7][11] ) );
  DFFX1 \regfile_reg[7][10]  ( .D(n422), .CLK(clk), .Q(\regfile[7][10] ) );
  DFFX1 \regfile_reg[7][9]  ( .D(n421), .CLK(clk), .Q(\regfile[7][9] ) );
  DFFX1 \regfile_reg[7][8]  ( .D(n420), .CLK(clk), .Q(\regfile[7][8] ) );
  DFFX1 \regfile_reg[7][7]  ( .D(n419), .CLK(clk), .Q(\regfile[7][7] ) );
  DFFX1 \regfile_reg[7][6]  ( .D(n418), .CLK(clk), .Q(\regfile[7][6] ) );
  DFFX1 \regfile_reg[7][5]  ( .D(n417), .CLK(clk), .Q(\regfile[7][5] ) );
  DFFX1 \regfile_reg[7][4]  ( .D(n416), .CLK(clk), .Q(\regfile[7][4] ) );
  DFFX1 \regfile_reg[7][3]  ( .D(n415), .CLK(clk), .Q(\regfile[7][3] ) );
  DFFX1 \regfile_reg[7][2]  ( .D(n414), .CLK(clk), .Q(\regfile[7][2] ) );
  DFFX1 \regfile_reg[7][1]  ( .D(n413), .CLK(clk), .Q(\regfile[7][1] ) );
  DFFX1 \regfile_reg[7][0]  ( .D(n412), .CLK(clk), .Q(\regfile[7][0] ) );
  DFFX1 \regfile_reg[6][31]  ( .D(n411), .CLK(clk), .Q(\regfile[6][31] ) );
  DFFX1 \regfile_reg[6][30]  ( .D(n410), .CLK(clk), .Q(\regfile[6][30] ) );
  DFFX1 \regfile_reg[6][29]  ( .D(n409), .CLK(clk), .Q(\regfile[6][29] ) );
  DFFX1 \regfile_reg[6][28]  ( .D(n408), .CLK(clk), .Q(\regfile[6][28] ) );
  DFFX1 \regfile_reg[6][27]  ( .D(n407), .CLK(clk), .Q(\regfile[6][27] ) );
  DFFX1 \regfile_reg[6][26]  ( .D(n406), .CLK(clk), .Q(\regfile[6][26] ) );
  DFFX1 \regfile_reg[6][25]  ( .D(n405), .CLK(clk), .Q(\regfile[6][25] ) );
  DFFX1 \regfile_reg[6][24]  ( .D(n404), .CLK(clk), .Q(\regfile[6][24] ) );
  DFFX1 \regfile_reg[6][23]  ( .D(n403), .CLK(clk), .Q(\regfile[6][23] ) );
  DFFX1 \regfile_reg[6][22]  ( .D(n402), .CLK(clk), .Q(\regfile[6][22] ) );
  DFFX1 \regfile_reg[6][21]  ( .D(n401), .CLK(clk), .Q(\regfile[6][21] ) );
  DFFX1 \regfile_reg[6][20]  ( .D(n400), .CLK(clk), .Q(\regfile[6][20] ) );
  DFFX1 \regfile_reg[6][19]  ( .D(n399), .CLK(clk), .Q(\regfile[6][19] ) );
  DFFX1 \regfile_reg[6][18]  ( .D(n398), .CLK(clk), .Q(\regfile[6][18] ) );
  DFFX1 \regfile_reg[6][17]  ( .D(n397), .CLK(clk), .Q(\regfile[6][17] ) );
  DFFX1 \regfile_reg[6][16]  ( .D(n396), .CLK(clk), .Q(\regfile[6][16] ) );
  DFFX1 \regfile_reg[6][15]  ( .D(n395), .CLK(clk), .Q(\regfile[6][15] ) );
  DFFX1 \regfile_reg[6][14]  ( .D(n394), .CLK(clk), .Q(\regfile[6][14] ) );
  DFFX1 \regfile_reg[6][13]  ( .D(n393), .CLK(clk), .Q(\regfile[6][13] ) );
  DFFX1 \regfile_reg[6][12]  ( .D(n392), .CLK(clk), .Q(\regfile[6][12] ) );
  DFFX1 \regfile_reg[6][11]  ( .D(n391), .CLK(clk), .Q(\regfile[6][11] ) );
  DFFX1 \regfile_reg[6][10]  ( .D(n390), .CLK(clk), .Q(\regfile[6][10] ) );
  DFFX1 \regfile_reg[6][9]  ( .D(n389), .CLK(clk), .Q(\regfile[6][9] ) );
  DFFX1 \regfile_reg[6][8]  ( .D(n388), .CLK(clk), .Q(\regfile[6][8] ) );
  DFFX1 \regfile_reg[6][7]  ( .D(n387), .CLK(clk), .Q(\regfile[6][7] ) );
  DFFX1 \regfile_reg[6][6]  ( .D(n386), .CLK(clk), .Q(\regfile[6][6] ) );
  DFFX1 \regfile_reg[6][5]  ( .D(n385), .CLK(clk), .Q(\regfile[6][5] ) );
  DFFX1 \regfile_reg[6][4]  ( .D(n384), .CLK(clk), .Q(\regfile[6][4] ) );
  DFFX1 \regfile_reg[6][3]  ( .D(n383), .CLK(clk), .Q(\regfile[6][3] ) );
  DFFX1 \regfile_reg[6][2]  ( .D(n382), .CLK(clk), .Q(\regfile[6][2] ) );
  DFFX1 \regfile_reg[6][1]  ( .D(n381), .CLK(clk), .Q(\regfile[6][1] ) );
  DFFX1 \regfile_reg[6][0]  ( .D(n380), .CLK(clk), .Q(\regfile[6][0] ) );
  DFFX1 \regfile_reg[5][31]  ( .D(n379), .CLK(clk), .Q(\regfile[5][31] ) );
  DFFX1 \regfile_reg[5][30]  ( .D(n378), .CLK(clk), .Q(\regfile[5][30] ) );
  DFFX1 \regfile_reg[5][29]  ( .D(n377), .CLK(clk), .Q(\regfile[5][29] ) );
  DFFX1 \regfile_reg[5][28]  ( .D(n376), .CLK(clk), .Q(\regfile[5][28] ) );
  DFFX1 \regfile_reg[5][27]  ( .D(n375), .CLK(clk), .Q(\regfile[5][27] ) );
  DFFX1 \regfile_reg[5][26]  ( .D(n374), .CLK(clk), .Q(\regfile[5][26] ) );
  DFFX1 \regfile_reg[5][25]  ( .D(n373), .CLK(clk), .Q(\regfile[5][25] ) );
  DFFX1 \regfile_reg[5][24]  ( .D(n372), .CLK(clk), .Q(\regfile[5][24] ) );
  DFFX1 \regfile_reg[5][23]  ( .D(n371), .CLK(clk), .Q(\regfile[5][23] ) );
  DFFX1 \regfile_reg[5][22]  ( .D(n370), .CLK(clk), .Q(\regfile[5][22] ) );
  DFFX1 \regfile_reg[5][21]  ( .D(n369), .CLK(clk), .Q(\regfile[5][21] ) );
  DFFX1 \regfile_reg[5][20]  ( .D(n368), .CLK(clk), .Q(\regfile[5][20] ) );
  DFFX1 \regfile_reg[5][19]  ( .D(n367), .CLK(clk), .Q(\regfile[5][19] ) );
  DFFX1 \regfile_reg[5][18]  ( .D(n366), .CLK(clk), .Q(\regfile[5][18] ) );
  DFFX1 \regfile_reg[5][17]  ( .D(n365), .CLK(clk), .Q(\regfile[5][17] ) );
  DFFX1 \regfile_reg[5][16]  ( .D(n364), .CLK(clk), .Q(\regfile[5][16] ) );
  DFFX1 \regfile_reg[5][15]  ( .D(n363), .CLK(clk), .Q(\regfile[5][15] ) );
  DFFX1 \regfile_reg[5][14]  ( .D(n362), .CLK(clk), .Q(\regfile[5][14] ) );
  DFFX1 \regfile_reg[5][13]  ( .D(n361), .CLK(clk), .Q(\regfile[5][13] ) );
  DFFX1 \regfile_reg[5][12]  ( .D(n360), .CLK(clk), .Q(\regfile[5][12] ) );
  DFFX1 \regfile_reg[5][11]  ( .D(n359), .CLK(clk), .Q(\regfile[5][11] ) );
  DFFX1 \regfile_reg[5][10]  ( .D(n358), .CLK(clk), .Q(\regfile[5][10] ) );
  DFFX1 \regfile_reg[5][9]  ( .D(n357), .CLK(clk), .Q(\regfile[5][9] ) );
  DFFX1 \regfile_reg[5][8]  ( .D(n356), .CLK(clk), .Q(\regfile[5][8] ) );
  DFFX1 \regfile_reg[5][7]  ( .D(n355), .CLK(clk), .Q(\regfile[5][7] ) );
  DFFX1 \regfile_reg[5][6]  ( .D(n354), .CLK(clk), .Q(\regfile[5][6] ) );
  DFFX1 \regfile_reg[5][5]  ( .D(n353), .CLK(clk), .Q(\regfile[5][5] ) );
  DFFX1 \regfile_reg[5][4]  ( .D(n352), .CLK(clk), .Q(\regfile[5][4] ) );
  DFFX1 \regfile_reg[5][3]  ( .D(n351), .CLK(clk), .Q(\regfile[5][3] ) );
  DFFX1 \regfile_reg[5][2]  ( .D(n350), .CLK(clk), .Q(\regfile[5][2] ) );
  DFFX1 \regfile_reg[5][1]  ( .D(n349), .CLK(clk), .Q(\regfile[5][1] ) );
  DFFX1 \regfile_reg[5][0]  ( .D(n348), .CLK(clk), .Q(\regfile[5][0] ) );
  DFFX1 \regfile_reg[4][31]  ( .D(n347), .CLK(clk), .Q(\regfile[4][31] ) );
  DFFX1 \regfile_reg[4][30]  ( .D(n346), .CLK(clk), .Q(\regfile[4][30] ) );
  DFFX1 \regfile_reg[4][29]  ( .D(n345), .CLK(clk), .Q(\regfile[4][29] ) );
  DFFX1 \regfile_reg[4][28]  ( .D(n344), .CLK(clk), .Q(\regfile[4][28] ) );
  DFFX1 \regfile_reg[4][27]  ( .D(n343), .CLK(clk), .Q(\regfile[4][27] ) );
  DFFX1 \regfile_reg[4][26]  ( .D(n342), .CLK(clk), .Q(\regfile[4][26] ) );
  DFFX1 \regfile_reg[4][25]  ( .D(n341), .CLK(clk), .Q(\regfile[4][25] ) );
  DFFX1 \regfile_reg[4][24]  ( .D(n340), .CLK(clk), .Q(\regfile[4][24] ) );
  DFFX1 \regfile_reg[4][23]  ( .D(n339), .CLK(clk), .Q(\regfile[4][23] ) );
  DFFX1 \regfile_reg[4][22]  ( .D(n338), .CLK(clk), .Q(\regfile[4][22] ) );
  DFFX1 \regfile_reg[4][21]  ( .D(n337), .CLK(clk), .Q(\regfile[4][21] ) );
  DFFX1 \regfile_reg[4][20]  ( .D(n336), .CLK(clk), .Q(\regfile[4][20] ) );
  DFFX1 \regfile_reg[4][19]  ( .D(n335), .CLK(clk), .Q(\regfile[4][19] ) );
  DFFX1 \regfile_reg[4][18]  ( .D(n334), .CLK(clk), .Q(\regfile[4][18] ) );
  DFFX1 \regfile_reg[4][17]  ( .D(n333), .CLK(clk), .Q(\regfile[4][17] ) );
  DFFX1 \regfile_reg[4][16]  ( .D(n332), .CLK(clk), .Q(\regfile[4][16] ) );
  DFFX1 \regfile_reg[4][15]  ( .D(n331), .CLK(clk), .Q(\regfile[4][15] ) );
  DFFX1 \regfile_reg[4][14]  ( .D(n330), .CLK(clk), .Q(\regfile[4][14] ) );
  DFFX1 \regfile_reg[4][13]  ( .D(n329), .CLK(clk), .Q(\regfile[4][13] ) );
  DFFX1 \regfile_reg[4][12]  ( .D(n328), .CLK(clk), .Q(\regfile[4][12] ) );
  DFFX1 \regfile_reg[4][11]  ( .D(n327), .CLK(clk), .Q(\regfile[4][11] ) );
  DFFX1 \regfile_reg[4][10]  ( .D(n326), .CLK(clk), .Q(\regfile[4][10] ) );
  DFFX1 \regfile_reg[4][9]  ( .D(n325), .CLK(clk), .Q(\regfile[4][9] ) );
  DFFX1 \regfile_reg[4][8]  ( .D(n324), .CLK(clk), .Q(\regfile[4][8] ) );
  DFFX1 \regfile_reg[4][7]  ( .D(n323), .CLK(clk), .Q(\regfile[4][7] ) );
  DFFX1 \regfile_reg[4][6]  ( .D(n322), .CLK(clk), .Q(\regfile[4][6] ) );
  DFFX1 \regfile_reg[4][5]  ( .D(n321), .CLK(clk), .Q(\regfile[4][5] ) );
  DFFX1 \regfile_reg[4][4]  ( .D(n320), .CLK(clk), .Q(\regfile[4][4] ) );
  DFFX1 \regfile_reg[4][3]  ( .D(n319), .CLK(clk), .Q(\regfile[4][3] ) );
  DFFX1 \regfile_reg[4][2]  ( .D(n318), .CLK(clk), .Q(\regfile[4][2] ) );
  DFFX1 \regfile_reg[4][1]  ( .D(n317), .CLK(clk), .Q(\regfile[4][1] ) );
  DFFX1 \regfile_reg[4][0]  ( .D(n316), .CLK(clk), .Q(\regfile[4][0] ) );
  DFFX1 \regfile_reg[3][31]  ( .D(n315), .CLK(clk), .Q(\regfile[3][31] ) );
  DFFX1 \regfile_reg[3][30]  ( .D(n314), .CLK(clk), .Q(\regfile[3][30] ) );
  DFFX1 \regfile_reg[3][29]  ( .D(n313), .CLK(clk), .Q(\regfile[3][29] ) );
  DFFX1 \regfile_reg[3][28]  ( .D(n312), .CLK(clk), .Q(\regfile[3][28] ) );
  DFFX1 \regfile_reg[3][27]  ( .D(n311), .CLK(clk), .Q(\regfile[3][27] ) );
  DFFX1 \regfile_reg[3][26]  ( .D(n310), .CLK(clk), .Q(\regfile[3][26] ) );
  DFFX1 \regfile_reg[3][25]  ( .D(n309), .CLK(clk), .Q(\regfile[3][25] ) );
  DFFX1 \regfile_reg[3][24]  ( .D(n308), .CLK(clk), .Q(\regfile[3][24] ) );
  DFFX1 \regfile_reg[3][23]  ( .D(n307), .CLK(clk), .Q(\regfile[3][23] ) );
  DFFX1 \regfile_reg[3][22]  ( .D(n306), .CLK(clk), .Q(\regfile[3][22] ) );
  DFFX1 \regfile_reg[3][21]  ( .D(n305), .CLK(clk), .Q(\regfile[3][21] ) );
  DFFX1 \regfile_reg[3][20]  ( .D(n304), .CLK(clk), .Q(\regfile[3][20] ) );
  DFFX1 \regfile_reg[3][19]  ( .D(n303), .CLK(clk), .Q(\regfile[3][19] ) );
  DFFX1 \regfile_reg[3][18]  ( .D(n302), .CLK(clk), .Q(\regfile[3][18] ) );
  DFFX1 \regfile_reg[3][17]  ( .D(n301), .CLK(clk), .Q(\regfile[3][17] ) );
  DFFX1 \regfile_reg[3][16]  ( .D(n300), .CLK(clk), .Q(\regfile[3][16] ) );
  DFFX1 \regfile_reg[3][15]  ( .D(n299), .CLK(clk), .Q(\regfile[3][15] ) );
  DFFX1 \regfile_reg[3][14]  ( .D(n298), .CLK(clk), .Q(\regfile[3][14] ) );
  DFFX1 \regfile_reg[3][13]  ( .D(n297), .CLK(clk), .Q(\regfile[3][13] ) );
  DFFX1 \regfile_reg[3][12]  ( .D(n296), .CLK(clk), .Q(\regfile[3][12] ) );
  DFFX1 \regfile_reg[3][11]  ( .D(n295), .CLK(clk), .Q(\regfile[3][11] ) );
  DFFX1 \regfile_reg[3][10]  ( .D(n294), .CLK(clk), .Q(\regfile[3][10] ) );
  DFFX1 \regfile_reg[3][9]  ( .D(n293), .CLK(clk), .Q(\regfile[3][9] ) );
  DFFX1 \regfile_reg[3][8]  ( .D(n292), .CLK(clk), .Q(\regfile[3][8] ) );
  DFFX1 \regfile_reg[3][7]  ( .D(n291), .CLK(clk), .Q(\regfile[3][7] ) );
  DFFX1 \regfile_reg[3][6]  ( .D(n290), .CLK(clk), .Q(\regfile[3][6] ) );
  DFFX1 \regfile_reg[3][5]  ( .D(n289), .CLK(clk), .Q(\regfile[3][5] ) );
  DFFX1 \regfile_reg[3][4]  ( .D(n288), .CLK(clk), .Q(\regfile[3][4] ) );
  DFFX1 \regfile_reg[3][3]  ( .D(n287), .CLK(clk), .Q(\regfile[3][3] ) );
  DFFX1 \regfile_reg[3][2]  ( .D(n286), .CLK(clk), .Q(\regfile[3][2] ) );
  DFFX1 \regfile_reg[3][1]  ( .D(n285), .CLK(clk), .Q(\regfile[3][1] ) );
  DFFX1 \regfile_reg[3][0]  ( .D(n284), .CLK(clk), .Q(\regfile[3][0] ) );
  DFFX1 \regfile_reg[2][31]  ( .D(n283), .CLK(clk), .Q(\regfile[2][31] ) );
  DFFX1 \regfile_reg[2][30]  ( .D(n282), .CLK(clk), .Q(\regfile[2][30] ) );
  DFFX1 \regfile_reg[2][29]  ( .D(n281), .CLK(clk), .Q(\regfile[2][29] ) );
  DFFX1 \regfile_reg[2][28]  ( .D(n280), .CLK(clk), .Q(\regfile[2][28] ) );
  DFFX1 \regfile_reg[2][27]  ( .D(n279), .CLK(clk), .Q(\regfile[2][27] ) );
  DFFX1 \regfile_reg[2][26]  ( .D(n278), .CLK(clk), .Q(\regfile[2][26] ) );
  DFFX1 \regfile_reg[2][25]  ( .D(n277), .CLK(clk), .Q(\regfile[2][25] ) );
  DFFX1 \regfile_reg[2][24]  ( .D(n276), .CLK(clk), .Q(\regfile[2][24] ) );
  DFFX1 \regfile_reg[2][23]  ( .D(n275), .CLK(clk), .Q(\regfile[2][23] ) );
  DFFX1 \regfile_reg[2][22]  ( .D(n274), .CLK(clk), .Q(\regfile[2][22] ) );
  DFFX1 \regfile_reg[2][21]  ( .D(n273), .CLK(clk), .Q(\regfile[2][21] ) );
  DFFX1 \regfile_reg[2][20]  ( .D(n272), .CLK(clk), .Q(\regfile[2][20] ) );
  DFFX1 \regfile_reg[2][19]  ( .D(n271), .CLK(clk), .Q(\regfile[2][19] ) );
  DFFX1 \regfile_reg[2][18]  ( .D(n270), .CLK(clk), .Q(\regfile[2][18] ) );
  DFFX1 \regfile_reg[2][17]  ( .D(n269), .CLK(clk), .Q(\regfile[2][17] ) );
  DFFX1 \regfile_reg[2][16]  ( .D(n268), .CLK(clk), .Q(\regfile[2][16] ) );
  DFFX1 \regfile_reg[2][15]  ( .D(n267), .CLK(clk), .Q(\regfile[2][15] ) );
  DFFX1 \regfile_reg[2][14]  ( .D(n266), .CLK(clk), .Q(\regfile[2][14] ) );
  DFFX1 \regfile_reg[2][13]  ( .D(n265), .CLK(clk), .Q(\regfile[2][13] ) );
  DFFX1 \regfile_reg[2][12]  ( .D(n264), .CLK(clk), .Q(\regfile[2][12] ) );
  DFFX1 \regfile_reg[2][11]  ( .D(n263), .CLK(clk), .Q(\regfile[2][11] ) );
  DFFX1 \regfile_reg[2][10]  ( .D(n262), .CLK(clk), .Q(\regfile[2][10] ) );
  DFFX1 \regfile_reg[2][9]  ( .D(n261), .CLK(clk), .Q(\regfile[2][9] ) );
  DFFX1 \regfile_reg[2][8]  ( .D(n260), .CLK(clk), .Q(\regfile[2][8] ) );
  DFFX1 \regfile_reg[2][7]  ( .D(n259), .CLK(clk), .Q(\regfile[2][7] ) );
  DFFX1 \regfile_reg[2][6]  ( .D(n258), .CLK(clk), .Q(\regfile[2][6] ) );
  DFFX1 \regfile_reg[2][5]  ( .D(n257), .CLK(clk), .Q(\regfile[2][5] ) );
  DFFX1 \regfile_reg[2][4]  ( .D(n256), .CLK(clk), .Q(\regfile[2][4] ) );
  DFFX1 \regfile_reg[2][3]  ( .D(n255), .CLK(clk), .Q(\regfile[2][3] ) );
  DFFX1 \regfile_reg[2][2]  ( .D(n254), .CLK(clk), .Q(\regfile[2][2] ) );
  DFFX1 \regfile_reg[2][1]  ( .D(n253), .CLK(clk), .Q(\regfile[2][1] ) );
  DFFX1 \regfile_reg[2][0]  ( .D(n252), .CLK(clk), .Q(\regfile[2][0] ) );
  DFFX1 \regfile_reg[1][31]  ( .D(n251), .CLK(clk), .Q(\regfile[1][31] ) );
  DFFX1 \regfile_reg[1][30]  ( .D(n250), .CLK(clk), .Q(\regfile[1][30] ) );
  DFFX1 \regfile_reg[1][29]  ( .D(n249), .CLK(clk), .Q(\regfile[1][29] ) );
  DFFX1 \regfile_reg[1][28]  ( .D(n248), .CLK(clk), .Q(\regfile[1][28] ) );
  DFFX1 \regfile_reg[1][27]  ( .D(n247), .CLK(clk), .Q(\regfile[1][27] ) );
  DFFX1 \regfile_reg[1][26]  ( .D(n246), .CLK(clk), .Q(\regfile[1][26] ) );
  DFFX1 \regfile_reg[1][25]  ( .D(n245), .CLK(clk), .Q(\regfile[1][25] ) );
  DFFX1 \regfile_reg[1][24]  ( .D(n244), .CLK(clk), .Q(\regfile[1][24] ) );
  DFFX1 \regfile_reg[1][23]  ( .D(n243), .CLK(clk), .Q(\regfile[1][23] ) );
  DFFX1 \regfile_reg[1][22]  ( .D(n242), .CLK(clk), .Q(\regfile[1][22] ) );
  DFFX1 \regfile_reg[1][21]  ( .D(n241), .CLK(clk), .Q(\regfile[1][21] ) );
  DFFX1 \regfile_reg[1][20]  ( .D(n240), .CLK(clk), .Q(\regfile[1][20] ) );
  DFFX1 \regfile_reg[1][19]  ( .D(n239), .CLK(clk), .Q(\regfile[1][19] ) );
  DFFX1 \regfile_reg[1][18]  ( .D(n238), .CLK(clk), .Q(\regfile[1][18] ) );
  DFFX1 \regfile_reg[1][17]  ( .D(n237), .CLK(clk), .Q(\regfile[1][17] ) );
  DFFX1 \regfile_reg[1][16]  ( .D(n236), .CLK(clk), .Q(\regfile[1][16] ) );
  DFFX1 \regfile_reg[1][15]  ( .D(n235), .CLK(clk), .Q(\regfile[1][15] ) );
  DFFX1 \regfile_reg[1][14]  ( .D(n234), .CLK(clk), .Q(\regfile[1][14] ) );
  DFFX1 \regfile_reg[1][13]  ( .D(n233), .CLK(clk), .Q(\regfile[1][13] ) );
  DFFX1 \regfile_reg[1][12]  ( .D(n232), .CLK(clk), .Q(\regfile[1][12] ) );
  DFFX1 \regfile_reg[1][11]  ( .D(n231), .CLK(clk), .Q(\regfile[1][11] ) );
  DFFX1 \regfile_reg[1][10]  ( .D(n230), .CLK(clk), .Q(\regfile[1][10] ) );
  DFFX1 \regfile_reg[1][9]  ( .D(n229), .CLK(clk), .Q(\regfile[1][9] ) );
  DFFX1 \regfile_reg[1][8]  ( .D(n228), .CLK(clk), .Q(\regfile[1][8] ) );
  DFFX1 \regfile_reg[1][7]  ( .D(n227), .CLK(clk), .Q(\regfile[1][7] ) );
  DFFX1 \regfile_reg[1][6]  ( .D(n226), .CLK(clk), .Q(\regfile[1][6] ) );
  DFFX1 \regfile_reg[1][5]  ( .D(n225), .CLK(clk), .Q(\regfile[1][5] ) );
  DFFX1 \regfile_reg[1][4]  ( .D(n224), .CLK(clk), .Q(\regfile[1][4] ) );
  DFFX1 \regfile_reg[1][3]  ( .D(n223), .CLK(clk), .Q(\regfile[1][3] ) );
  DFFX1 \regfile_reg[1][2]  ( .D(n222), .CLK(clk), .Q(\regfile[1][2] ) );
  DFFX1 \regfile_reg[1][1]  ( .D(n221), .CLK(clk), .Q(\regfile[1][1] ) );
  DFFX1 \regfile_reg[1][0]  ( .D(n220), .CLK(clk), .Q(\regfile[1][0] ) );
  DFFX1 \regfile_reg[0][31]  ( .D(n219), .CLK(clk), .Q(\regfile[0][31] ) );
  DFFX1 \regfile_reg[0][30]  ( .D(n218), .CLK(clk), .Q(\regfile[0][30] ) );
  DFFX1 \regfile_reg[0][29]  ( .D(n217), .CLK(clk), .Q(\regfile[0][29] ) );
  DFFX1 \regfile_reg[0][28]  ( .D(n216), .CLK(clk), .Q(\regfile[0][28] ) );
  DFFX1 \regfile_reg[0][27]  ( .D(n215), .CLK(clk), .Q(\regfile[0][27] ) );
  DFFX1 \regfile_reg[0][26]  ( .D(n214), .CLK(clk), .Q(\regfile[0][26] ) );
  DFFX1 \regfile_reg[0][25]  ( .D(n213), .CLK(clk), .Q(\regfile[0][25] ) );
  DFFX1 \regfile_reg[0][24]  ( .D(n212), .CLK(clk), .Q(\regfile[0][24] ) );
  DFFX1 \regfile_reg[0][23]  ( .D(n211), .CLK(clk), .Q(\regfile[0][23] ) );
  DFFX1 \regfile_reg[0][22]  ( .D(n210), .CLK(clk), .Q(\regfile[0][22] ) );
  DFFX1 \regfile_reg[0][21]  ( .D(n209), .CLK(clk), .Q(\regfile[0][21] ) );
  DFFX1 \regfile_reg[0][20]  ( .D(n208), .CLK(clk), .Q(\regfile[0][20] ) );
  DFFX1 \regfile_reg[0][19]  ( .D(n207), .CLK(clk), .Q(\regfile[0][19] ) );
  DFFX1 \regfile_reg[0][18]  ( .D(n206), .CLK(clk), .Q(\regfile[0][18] ) );
  DFFX1 \regfile_reg[0][17]  ( .D(n205), .CLK(clk), .Q(\regfile[0][17] ) );
  DFFX1 \regfile_reg[0][16]  ( .D(n204), .CLK(clk), .Q(\regfile[0][16] ) );
  DFFX1 \regfile_reg[0][15]  ( .D(n203), .CLK(clk), .Q(\regfile[0][15] ) );
  DFFX1 \regfile_reg[0][14]  ( .D(n202), .CLK(clk), .Q(\regfile[0][14] ) );
  DFFX1 \regfile_reg[0][13]  ( .D(n201), .CLK(clk), .Q(\regfile[0][13] ) );
  DFFX1 \regfile_reg[0][12]  ( .D(n200), .CLK(clk), .Q(\regfile[0][12] ) );
  DFFX1 \regfile_reg[0][11]  ( .D(n199), .CLK(clk), .Q(\regfile[0][11] ) );
  DFFX1 \regfile_reg[0][10]  ( .D(n198), .CLK(clk), .Q(\regfile[0][10] ) );
  DFFX1 \regfile_reg[0][9]  ( .D(n197), .CLK(clk), .Q(\regfile[0][9] ) );
  DFFX1 \regfile_reg[0][8]  ( .D(n196), .CLK(clk), .Q(\regfile[0][8] ) );
  DFFX1 \regfile_reg[0][7]  ( .D(n195), .CLK(clk), .Q(\regfile[0][7] ) );
  DFFX1 \regfile_reg[0][6]  ( .D(n194), .CLK(clk), .Q(\regfile[0][6] ) );
  DFFX1 \regfile_reg[0][5]  ( .D(n193), .CLK(clk), .Q(\regfile[0][5] ) );
  DFFX1 \regfile_reg[0][4]  ( .D(n192), .CLK(clk), .Q(\regfile[0][4] ) );
  DFFX1 \regfile_reg[0][3]  ( .D(n191), .CLK(clk), .Q(\regfile[0][3] ) );
  DFFX1 \regfile_reg[0][2]  ( .D(n190), .CLK(clk), .Q(\regfile[0][2] ) );
  DFFX1 \regfile_reg[0][1]  ( .D(n189), .CLK(clk), .Q(\regfile[0][1] ) );
  DFFX1 \regfile_reg[0][0]  ( .D(n188), .CLK(clk), .Q(\regfile[0][0] ) );
  AO22X1 U3 ( .IN1(n1169), .IN2(N299), .IN3(\regfile[9][9] ), .IN4(n1164), .Q(
        n485) );
  AO22X1 U4 ( .IN1(n1169), .IN2(N298), .IN3(\regfile[9][8] ), .IN4(n1164), .Q(
        n484) );
  AO22X1 U5 ( .IN1(n1169), .IN2(N297), .IN3(\regfile[9][7] ), .IN4(n1164), .Q(
        n483) );
  AO22X1 U6 ( .IN1(n1169), .IN2(N296), .IN3(\regfile[9][6] ), .IN4(n1164), .Q(
        n482) );
  AO22X1 U11 ( .IN1(n1169), .IN2(N295), .IN3(\regfile[9][5] ), .IN4(n1164), 
        .Q(n481) );
  AO22X1 U12 ( .IN1(n1169), .IN2(N294), .IN3(\regfile[9][4] ), .IN4(n1164), 
        .Q(n480) );
  AO22X1 U13 ( .IN1(n1169), .IN2(N293), .IN3(\regfile[9][3] ), .IN4(n1164), 
        .Q(n479) );
  AO22X1 U14 ( .IN1(n1168), .IN2(N321), .IN3(\regfile[9][31] ), .IN4(n1164), 
        .Q(n507) );
  AO22X1 U15 ( .IN1(n1168), .IN2(N320), .IN3(\regfile[9][30] ), .IN4(n1163), 
        .Q(n506) );
  AO22X1 U16 ( .IN1(n1168), .IN2(N292), .IN3(\regfile[9][2] ), .IN4(n1163), 
        .Q(n478) );
  AO22X1 U17 ( .IN1(n1168), .IN2(N319), .IN3(\regfile[9][29] ), .IN4(n1163), 
        .Q(n505) );
  AO22X1 U18 ( .IN1(n1168), .IN2(N318), .IN3(\regfile[9][28] ), .IN4(n1163), 
        .Q(n504) );
  AO22X1 U19 ( .IN1(n1168), .IN2(N317), .IN3(\regfile[9][27] ), .IN4(n1163), 
        .Q(n503) );
  AO22X1 U20 ( .IN1(n1168), .IN2(N316), .IN3(\regfile[9][26] ), .IN4(n1163), 
        .Q(n502) );
  AO22X1 U21 ( .IN1(n1167), .IN2(N315), .IN3(\regfile[9][25] ), .IN4(n1163), 
        .Q(n501) );
  AO22X1 U22 ( .IN1(n1167), .IN2(N314), .IN3(\regfile[9][24] ), .IN4(n1163), 
        .Q(n500) );
  AO22X1 U23 ( .IN1(n1167), .IN2(N313), .IN3(\regfile[9][23] ), .IN4(n1163), 
        .Q(n499) );
  AO22X1 U24 ( .IN1(n1167), .IN2(N312), .IN3(\regfile[9][22] ), .IN4(n1163), 
        .Q(n498) );
  AO22X1 U25 ( .IN1(n1167), .IN2(N311), .IN3(\regfile[9][21] ), .IN4(n1163), 
        .Q(n497) );
  AO22X1 U26 ( .IN1(n1167), .IN2(N310), .IN3(\regfile[9][20] ), .IN4(n1163), 
        .Q(n496) );
  AO22X1 U27 ( .IN1(n1167), .IN2(N291), .IN3(\regfile[9][1] ), .IN4(n1162), 
        .Q(n477) );
  AO22X1 U28 ( .IN1(n1166), .IN2(N309), .IN3(\regfile[9][19] ), .IN4(n1162), 
        .Q(n495) );
  AO22X1 U29 ( .IN1(n1166), .IN2(N308), .IN3(\regfile[9][18] ), .IN4(n1162), 
        .Q(n494) );
  AO22X1 U30 ( .IN1(n1166), .IN2(N307), .IN3(\regfile[9][17] ), .IN4(n1162), 
        .Q(n493) );
  AO22X1 U31 ( .IN1(n1166), .IN2(N306), .IN3(\regfile[9][16] ), .IN4(n1162), 
        .Q(n492) );
  AO22X1 U32 ( .IN1(n1166), .IN2(N305), .IN3(\regfile[9][15] ), .IN4(n1162), 
        .Q(n491) );
  AO22X1 U33 ( .IN1(n1166), .IN2(N304), .IN3(\regfile[9][14] ), .IN4(n1162), 
        .Q(n490) );
  AO22X1 U34 ( .IN1(n1166), .IN2(N303), .IN3(\regfile[9][13] ), .IN4(n1162), 
        .Q(n489) );
  AO22X1 U35 ( .IN1(n1165), .IN2(N302), .IN3(\regfile[9][12] ), .IN4(n1162), 
        .Q(n488) );
  AO22X1 U36 ( .IN1(n1165), .IN2(N301), .IN3(\regfile[9][11] ), .IN4(n1162), 
        .Q(n487) );
  AO22X1 U37 ( .IN1(n1165), .IN2(N300), .IN3(\regfile[9][10] ), .IN4(n1162), 
        .Q(n486) );
  AO22X1 U38 ( .IN1(n1165), .IN2(N290), .IN3(\regfile[9][0] ), .IN4(n1162), 
        .Q(n476) );
  AO22X1 U41 ( .IN1(n1161), .IN2(N299), .IN3(\regfile[8][9] ), .IN4(n1156), 
        .Q(n453) );
  AO22X1 U42 ( .IN1(n1161), .IN2(N298), .IN3(\regfile[8][8] ), .IN4(n1156), 
        .Q(n452) );
  AO22X1 U43 ( .IN1(n1161), .IN2(N297), .IN3(\regfile[8][7] ), .IN4(n1156), 
        .Q(n451) );
  AO22X1 U44 ( .IN1(n1161), .IN2(N296), .IN3(\regfile[8][6] ), .IN4(n1156), 
        .Q(n450) );
  AO22X1 U45 ( .IN1(n1161), .IN2(N295), .IN3(\regfile[8][5] ), .IN4(n1156), 
        .Q(n449) );
  AO22X1 U46 ( .IN1(n1161), .IN2(N294), .IN3(\regfile[8][4] ), .IN4(n1156), 
        .Q(n448) );
  AO22X1 U47 ( .IN1(n1161), .IN2(N293), .IN3(\regfile[8][3] ), .IN4(n1156), 
        .Q(n447) );
  AO22X1 U48 ( .IN1(n1160), .IN2(N321), .IN3(\regfile[8][31] ), .IN4(n1156), 
        .Q(n475) );
  AO22X1 U49 ( .IN1(n1160), .IN2(N320), .IN3(\regfile[8][30] ), .IN4(n1155), 
        .Q(n474) );
  AO22X1 U50 ( .IN1(n1160), .IN2(N292), .IN3(\regfile[8][2] ), .IN4(n1155), 
        .Q(n446) );
  AO22X1 U51 ( .IN1(n1160), .IN2(N319), .IN3(\regfile[8][29] ), .IN4(n1155), 
        .Q(n473) );
  AO22X1 U52 ( .IN1(n1160), .IN2(N318), .IN3(\regfile[8][28] ), .IN4(n1155), 
        .Q(n472) );
  AO22X1 U53 ( .IN1(n1160), .IN2(N317), .IN3(\regfile[8][27] ), .IN4(n1155), 
        .Q(n471) );
  AO22X1 U54 ( .IN1(n1160), .IN2(N316), .IN3(\regfile[8][26] ), .IN4(n1155), 
        .Q(n470) );
  AO22X1 U55 ( .IN1(n1159), .IN2(N315), .IN3(\regfile[8][25] ), .IN4(n1155), 
        .Q(n469) );
  AO22X1 U56 ( .IN1(n1159), .IN2(N314), .IN3(\regfile[8][24] ), .IN4(n1155), 
        .Q(n468) );
  AO22X1 U57 ( .IN1(n1159), .IN2(N313), .IN3(\regfile[8][23] ), .IN4(n1155), 
        .Q(n467) );
  AO22X1 U58 ( .IN1(n1159), .IN2(N312), .IN3(\regfile[8][22] ), .IN4(n1155), 
        .Q(n466) );
  AO22X1 U59 ( .IN1(n1159), .IN2(N311), .IN3(\regfile[8][21] ), .IN4(n1155), 
        .Q(n465) );
  AO22X1 U60 ( .IN1(n1159), .IN2(N310), .IN3(\regfile[8][20] ), .IN4(n1155), 
        .Q(n464) );
  AO22X1 U61 ( .IN1(n1159), .IN2(N291), .IN3(\regfile[8][1] ), .IN4(n1154), 
        .Q(n445) );
  AO22X1 U62 ( .IN1(n1158), .IN2(N309), .IN3(\regfile[8][19] ), .IN4(n1154), 
        .Q(n463) );
  AO22X1 U63 ( .IN1(n1158), .IN2(N308), .IN3(\regfile[8][18] ), .IN4(n1154), 
        .Q(n462) );
  AO22X1 U64 ( .IN1(n1158), .IN2(N307), .IN3(\regfile[8][17] ), .IN4(n1154), 
        .Q(n461) );
  AO22X1 U65 ( .IN1(n1158), .IN2(N306), .IN3(\regfile[8][16] ), .IN4(n1154), 
        .Q(n460) );
  AO22X1 U66 ( .IN1(n1158), .IN2(N305), .IN3(\regfile[8][15] ), .IN4(n1154), 
        .Q(n459) );
  AO22X1 U67 ( .IN1(n1158), .IN2(N304), .IN3(\regfile[8][14] ), .IN4(n1154), 
        .Q(n458) );
  AO22X1 U68 ( .IN1(n1158), .IN2(N303), .IN3(\regfile[8][13] ), .IN4(n1154), 
        .Q(n457) );
  AO22X1 U69 ( .IN1(n1157), .IN2(N302), .IN3(\regfile[8][12] ), .IN4(n1154), 
        .Q(n456) );
  AO22X1 U70 ( .IN1(n1157), .IN2(N301), .IN3(\regfile[8][11] ), .IN4(n1154), 
        .Q(n455) );
  AO22X1 U71 ( .IN1(n1157), .IN2(N300), .IN3(\regfile[8][10] ), .IN4(n1154), 
        .Q(n454) );
  AO22X1 U72 ( .IN1(n1157), .IN2(N290), .IN3(\regfile[8][0] ), .IN4(n1154), 
        .Q(n444) );
  AO22X1 U75 ( .IN1(n1153), .IN2(N299), .IN3(\regfile[7][9] ), .IN4(n1148), 
        .Q(n421) );
  AO22X1 U76 ( .IN1(n1153), .IN2(N298), .IN3(\regfile[7][8] ), .IN4(n1148), 
        .Q(n420) );
  AO22X1 U77 ( .IN1(n1153), .IN2(N297), .IN3(\regfile[7][7] ), .IN4(n1148), 
        .Q(n419) );
  AO22X1 U78 ( .IN1(n1153), .IN2(N296), .IN3(\regfile[7][6] ), .IN4(n1148), 
        .Q(n418) );
  AO22X1 U79 ( .IN1(n1153), .IN2(N295), .IN3(\regfile[7][5] ), .IN4(n1148), 
        .Q(n417) );
  AO22X1 U80 ( .IN1(n1153), .IN2(N294), .IN3(\regfile[7][4] ), .IN4(n1148), 
        .Q(n416) );
  AO22X1 U81 ( .IN1(n1153), .IN2(N293), .IN3(\regfile[7][3] ), .IN4(n1148), 
        .Q(n415) );
  AO22X1 U82 ( .IN1(n1152), .IN2(N321), .IN3(\regfile[7][31] ), .IN4(n1148), 
        .Q(n443) );
  AO22X1 U83 ( .IN1(n1152), .IN2(N320), .IN3(\regfile[7][30] ), .IN4(n1147), 
        .Q(n442) );
  AO22X1 U84 ( .IN1(n1152), .IN2(N292), .IN3(\regfile[7][2] ), .IN4(n1147), 
        .Q(n414) );
  AO22X1 U85 ( .IN1(n1152), .IN2(N319), .IN3(\regfile[7][29] ), .IN4(n1147), 
        .Q(n441) );
  AO22X1 U86 ( .IN1(n1152), .IN2(N318), .IN3(\regfile[7][28] ), .IN4(n1147), 
        .Q(n440) );
  AO22X1 U87 ( .IN1(n1152), .IN2(N317), .IN3(\regfile[7][27] ), .IN4(n1147), 
        .Q(n439) );
  AO22X1 U88 ( .IN1(n1152), .IN2(N316), .IN3(\regfile[7][26] ), .IN4(n1147), 
        .Q(n438) );
  AO22X1 U89 ( .IN1(n1151), .IN2(N315), .IN3(\regfile[7][25] ), .IN4(n1147), 
        .Q(n437) );
  AO22X1 U90 ( .IN1(n1151), .IN2(N314), .IN3(\regfile[7][24] ), .IN4(n1147), 
        .Q(n436) );
  AO22X1 U91 ( .IN1(n1151), .IN2(N313), .IN3(\regfile[7][23] ), .IN4(n1147), 
        .Q(n435) );
  AO22X1 U92 ( .IN1(n1151), .IN2(N312), .IN3(\regfile[7][22] ), .IN4(n1147), 
        .Q(n434) );
  AO22X1 U93 ( .IN1(n1151), .IN2(N311), .IN3(\regfile[7][21] ), .IN4(n1147), 
        .Q(n433) );
  AO22X1 U94 ( .IN1(n1151), .IN2(N310), .IN3(\regfile[7][20] ), .IN4(n1147), 
        .Q(n432) );
  AO22X1 U95 ( .IN1(n1151), .IN2(N291), .IN3(\regfile[7][1] ), .IN4(n1146), 
        .Q(n413) );
  AO22X1 U96 ( .IN1(n1150), .IN2(N309), .IN3(\regfile[7][19] ), .IN4(n1146), 
        .Q(n431) );
  AO22X1 U97 ( .IN1(n1150), .IN2(N308), .IN3(\regfile[7][18] ), .IN4(n1146), 
        .Q(n430) );
  AO22X1 U98 ( .IN1(n1150), .IN2(N307), .IN3(\regfile[7][17] ), .IN4(n1146), 
        .Q(n429) );
  AO22X1 U99 ( .IN1(n1150), .IN2(N306), .IN3(\regfile[7][16] ), .IN4(n1146), 
        .Q(n428) );
  AO22X1 U100 ( .IN1(n1150), .IN2(N305), .IN3(\regfile[7][15] ), .IN4(n1146), 
        .Q(n427) );
  AO22X1 U101 ( .IN1(n1150), .IN2(N304), .IN3(\regfile[7][14] ), .IN4(n1146), 
        .Q(n426) );
  AO22X1 U102 ( .IN1(n1150), .IN2(N303), .IN3(\regfile[7][13] ), .IN4(n1146), 
        .Q(n425) );
  AO22X1 U103 ( .IN1(n1149), .IN2(N302), .IN3(\regfile[7][12] ), .IN4(n1146), 
        .Q(n424) );
  AO22X1 U104 ( .IN1(n1149), .IN2(N301), .IN3(\regfile[7][11] ), .IN4(n1146), 
        .Q(n423) );
  AO22X1 U105 ( .IN1(n1149), .IN2(N300), .IN3(\regfile[7][10] ), .IN4(n1146), 
        .Q(n422) );
  AO22X1 U106 ( .IN1(n1149), .IN2(N290), .IN3(\regfile[7][0] ), .IN4(n1146), 
        .Q(n412) );
  AO22X1 U109 ( .IN1(n1145), .IN2(N299), .IN3(\regfile[6][9] ), .IN4(n1140), 
        .Q(n389) );
  AO22X1 U110 ( .IN1(n1145), .IN2(N298), .IN3(\regfile[6][8] ), .IN4(n1140), 
        .Q(n388) );
  AO22X1 U111 ( .IN1(n1145), .IN2(N297), .IN3(\regfile[6][7] ), .IN4(n1140), 
        .Q(n387) );
  AO22X1 U112 ( .IN1(n1145), .IN2(N296), .IN3(\regfile[6][6] ), .IN4(n1140), 
        .Q(n386) );
  AO22X1 U113 ( .IN1(n1145), .IN2(N295), .IN3(\regfile[6][5] ), .IN4(n1140), 
        .Q(n385) );
  AO22X1 U114 ( .IN1(n1145), .IN2(N294), .IN3(\regfile[6][4] ), .IN4(n1140), 
        .Q(n384) );
  AO22X1 U115 ( .IN1(n1145), .IN2(N293), .IN3(\regfile[6][3] ), .IN4(n1140), 
        .Q(n383) );
  AO22X1 U116 ( .IN1(n1144), .IN2(N321), .IN3(\regfile[6][31] ), .IN4(n1140), 
        .Q(n411) );
  AO22X1 U117 ( .IN1(n1144), .IN2(N320), .IN3(\regfile[6][30] ), .IN4(n1139), 
        .Q(n410) );
  AO22X1 U118 ( .IN1(n1144), .IN2(N292), .IN3(\regfile[6][2] ), .IN4(n1139), 
        .Q(n382) );
  AO22X1 U119 ( .IN1(n1144), .IN2(N319), .IN3(\regfile[6][29] ), .IN4(n1139), 
        .Q(n409) );
  AO22X1 U120 ( .IN1(n1144), .IN2(N318), .IN3(\regfile[6][28] ), .IN4(n1139), 
        .Q(n408) );
  AO22X1 U121 ( .IN1(n1144), .IN2(N317), .IN3(\regfile[6][27] ), .IN4(n1139), 
        .Q(n407) );
  AO22X1 U122 ( .IN1(n1144), .IN2(N316), .IN3(\regfile[6][26] ), .IN4(n1139), 
        .Q(n406) );
  AO22X1 U123 ( .IN1(n1143), .IN2(N315), .IN3(\regfile[6][25] ), .IN4(n1139), 
        .Q(n405) );
  AO22X1 U124 ( .IN1(n1143), .IN2(N314), .IN3(\regfile[6][24] ), .IN4(n1139), 
        .Q(n404) );
  AO22X1 U125 ( .IN1(n1143), .IN2(N313), .IN3(\regfile[6][23] ), .IN4(n1139), 
        .Q(n403) );
  AO22X1 U126 ( .IN1(n1143), .IN2(N312), .IN3(\regfile[6][22] ), .IN4(n1139), 
        .Q(n402) );
  AO22X1 U127 ( .IN1(n1143), .IN2(N311), .IN3(\regfile[6][21] ), .IN4(n1139), 
        .Q(n401) );
  AO22X1 U128 ( .IN1(n1143), .IN2(N310), .IN3(\regfile[6][20] ), .IN4(n1139), 
        .Q(n400) );
  AO22X1 U129 ( .IN1(n1143), .IN2(N291), .IN3(\regfile[6][1] ), .IN4(n1138), 
        .Q(n381) );
  AO22X1 U130 ( .IN1(n1142), .IN2(N309), .IN3(\regfile[6][19] ), .IN4(n1138), 
        .Q(n399) );
  AO22X1 U131 ( .IN1(n1142), .IN2(N308), .IN3(\regfile[6][18] ), .IN4(n1138), 
        .Q(n398) );
  AO22X1 U132 ( .IN1(n1142), .IN2(N307), .IN3(\regfile[6][17] ), .IN4(n1138), 
        .Q(n397) );
  AO22X1 U133 ( .IN1(n1142), .IN2(N306), .IN3(\regfile[6][16] ), .IN4(n1138), 
        .Q(n396) );
  AO22X1 U134 ( .IN1(n1142), .IN2(N305), .IN3(\regfile[6][15] ), .IN4(n1138), 
        .Q(n395) );
  AO22X1 U135 ( .IN1(n1142), .IN2(N304), .IN3(\regfile[6][14] ), .IN4(n1138), 
        .Q(n394) );
  AO22X1 U136 ( .IN1(n1142), .IN2(N303), .IN3(\regfile[6][13] ), .IN4(n1138), 
        .Q(n393) );
  AO22X1 U137 ( .IN1(n1141), .IN2(N302), .IN3(\regfile[6][12] ), .IN4(n1138), 
        .Q(n392) );
  AO22X1 U138 ( .IN1(n1141), .IN2(N301), .IN3(\regfile[6][11] ), .IN4(n1138), 
        .Q(n391) );
  AO22X1 U139 ( .IN1(n1141), .IN2(N300), .IN3(\regfile[6][10] ), .IN4(n1138), 
        .Q(n390) );
  AO22X1 U140 ( .IN1(n1141), .IN2(N290), .IN3(\regfile[6][0] ), .IN4(n1138), 
        .Q(n380) );
  AO22X1 U143 ( .IN1(n1137), .IN2(N299), .IN3(\regfile[5][9] ), .IN4(n1132), 
        .Q(n357) );
  AO22X1 U144 ( .IN1(n1137), .IN2(N298), .IN3(\regfile[5][8] ), .IN4(n1132), 
        .Q(n356) );
  AO22X1 U145 ( .IN1(n1137), .IN2(N297), .IN3(\regfile[5][7] ), .IN4(n1132), 
        .Q(n355) );
  AO22X1 U146 ( .IN1(n1137), .IN2(N296), .IN3(\regfile[5][6] ), .IN4(n1132), 
        .Q(n354) );
  AO22X1 U147 ( .IN1(n1137), .IN2(N295), .IN3(\regfile[5][5] ), .IN4(n1132), 
        .Q(n353) );
  AO22X1 U148 ( .IN1(n1137), .IN2(N294), .IN3(\regfile[5][4] ), .IN4(n1132), 
        .Q(n352) );
  AO22X1 U149 ( .IN1(n1137), .IN2(N293), .IN3(\regfile[5][3] ), .IN4(n1132), 
        .Q(n351) );
  AO22X1 U150 ( .IN1(n1136), .IN2(N321), .IN3(\regfile[5][31] ), .IN4(n1132), 
        .Q(n379) );
  AO22X1 U151 ( .IN1(n1136), .IN2(N320), .IN3(\regfile[5][30] ), .IN4(n1131), 
        .Q(n378) );
  AO22X1 U152 ( .IN1(n1136), .IN2(N292), .IN3(\regfile[5][2] ), .IN4(n1131), 
        .Q(n350) );
  AO22X1 U153 ( .IN1(n1136), .IN2(N319), .IN3(\regfile[5][29] ), .IN4(n1131), 
        .Q(n377) );
  AO22X1 U154 ( .IN1(n1136), .IN2(N318), .IN3(\regfile[5][28] ), .IN4(n1131), 
        .Q(n376) );
  AO22X1 U155 ( .IN1(n1136), .IN2(N317), .IN3(\regfile[5][27] ), .IN4(n1131), 
        .Q(n375) );
  AO22X1 U156 ( .IN1(n1136), .IN2(N316), .IN3(\regfile[5][26] ), .IN4(n1131), 
        .Q(n374) );
  AO22X1 U157 ( .IN1(n1135), .IN2(N315), .IN3(\regfile[5][25] ), .IN4(n1131), 
        .Q(n373) );
  AO22X1 U158 ( .IN1(n1135), .IN2(N314), .IN3(\regfile[5][24] ), .IN4(n1131), 
        .Q(n372) );
  AO22X1 U159 ( .IN1(n1135), .IN2(N313), .IN3(\regfile[5][23] ), .IN4(n1131), 
        .Q(n371) );
  AO22X1 U160 ( .IN1(n1135), .IN2(N312), .IN3(\regfile[5][22] ), .IN4(n1131), 
        .Q(n370) );
  AO22X1 U161 ( .IN1(n1135), .IN2(N311), .IN3(\regfile[5][21] ), .IN4(n1131), 
        .Q(n369) );
  AO22X1 U162 ( .IN1(n1135), .IN2(N310), .IN3(\regfile[5][20] ), .IN4(n1131), 
        .Q(n368) );
  AO22X1 U163 ( .IN1(n1135), .IN2(N291), .IN3(\regfile[5][1] ), .IN4(n1130), 
        .Q(n349) );
  AO22X1 U164 ( .IN1(n1134), .IN2(N309), .IN3(\regfile[5][19] ), .IN4(n1130), 
        .Q(n367) );
  AO22X1 U165 ( .IN1(n1134), .IN2(N308), .IN3(\regfile[5][18] ), .IN4(n1130), 
        .Q(n366) );
  AO22X1 U166 ( .IN1(n1134), .IN2(N307), .IN3(\regfile[5][17] ), .IN4(n1130), 
        .Q(n365) );
  AO22X1 U167 ( .IN1(n1134), .IN2(N306), .IN3(\regfile[5][16] ), .IN4(n1130), 
        .Q(n364) );
  AO22X1 U168 ( .IN1(n1134), .IN2(N305), .IN3(\regfile[5][15] ), .IN4(n1130), 
        .Q(n363) );
  AO22X1 U169 ( .IN1(n1134), .IN2(N304), .IN3(\regfile[5][14] ), .IN4(n1130), 
        .Q(n362) );
  AO22X1 U170 ( .IN1(n1134), .IN2(N303), .IN3(\regfile[5][13] ), .IN4(n1130), 
        .Q(n361) );
  AO22X1 U171 ( .IN1(n1133), .IN2(N302), .IN3(\regfile[5][12] ), .IN4(n1130), 
        .Q(n360) );
  AO22X1 U172 ( .IN1(n1133), .IN2(N301), .IN3(\regfile[5][11] ), .IN4(n1130), 
        .Q(n359) );
  AO22X1 U173 ( .IN1(n1133), .IN2(N300), .IN3(\regfile[5][10] ), .IN4(n1130), 
        .Q(n358) );
  AO22X1 U174 ( .IN1(n1133), .IN2(N290), .IN3(\regfile[5][0] ), .IN4(n1130), 
        .Q(n348) );
  AO22X1 U177 ( .IN1(n1129), .IN2(N299), .IN3(\regfile[4][9] ), .IN4(n1124), 
        .Q(n325) );
  AO22X1 U178 ( .IN1(n1129), .IN2(N298), .IN3(\regfile[4][8] ), .IN4(n1124), 
        .Q(n324) );
  AO22X1 U179 ( .IN1(n1129), .IN2(N297), .IN3(\regfile[4][7] ), .IN4(n1124), 
        .Q(n323) );
  AO22X1 U180 ( .IN1(n1129), .IN2(N296), .IN3(\regfile[4][6] ), .IN4(n1124), 
        .Q(n322) );
  AO22X1 U181 ( .IN1(n1129), .IN2(N295), .IN3(\regfile[4][5] ), .IN4(n1124), 
        .Q(n321) );
  AO22X1 U182 ( .IN1(n1129), .IN2(N294), .IN3(\regfile[4][4] ), .IN4(n1124), 
        .Q(n320) );
  AO22X1 U183 ( .IN1(n1129), .IN2(N293), .IN3(\regfile[4][3] ), .IN4(n1124), 
        .Q(n319) );
  AO22X1 U184 ( .IN1(n1128), .IN2(N321), .IN3(\regfile[4][31] ), .IN4(n1124), 
        .Q(n347) );
  AO22X1 U185 ( .IN1(n1128), .IN2(N320), .IN3(\regfile[4][30] ), .IN4(n1123), 
        .Q(n346) );
  AO22X1 U186 ( .IN1(n1128), .IN2(N292), .IN3(\regfile[4][2] ), .IN4(n1123), 
        .Q(n318) );
  AO22X1 U187 ( .IN1(n1128), .IN2(N319), .IN3(\regfile[4][29] ), .IN4(n1123), 
        .Q(n345) );
  AO22X1 U188 ( .IN1(n1128), .IN2(N318), .IN3(\regfile[4][28] ), .IN4(n1123), 
        .Q(n344) );
  AO22X1 U189 ( .IN1(n1128), .IN2(N317), .IN3(\regfile[4][27] ), .IN4(n1123), 
        .Q(n343) );
  AO22X1 U190 ( .IN1(n1128), .IN2(N316), .IN3(\regfile[4][26] ), .IN4(n1123), 
        .Q(n342) );
  AO22X1 U191 ( .IN1(n1127), .IN2(N315), .IN3(\regfile[4][25] ), .IN4(n1123), 
        .Q(n341) );
  AO22X1 U192 ( .IN1(n1127), .IN2(N314), .IN3(\regfile[4][24] ), .IN4(n1123), 
        .Q(n340) );
  AO22X1 U193 ( .IN1(n1127), .IN2(N313), .IN3(\regfile[4][23] ), .IN4(n1123), 
        .Q(n339) );
  AO22X1 U194 ( .IN1(n1127), .IN2(N312), .IN3(\regfile[4][22] ), .IN4(n1123), 
        .Q(n338) );
  AO22X1 U195 ( .IN1(n1127), .IN2(N311), .IN3(\regfile[4][21] ), .IN4(n1123), 
        .Q(n337) );
  AO22X1 U196 ( .IN1(n1127), .IN2(N310), .IN3(\regfile[4][20] ), .IN4(n1123), 
        .Q(n336) );
  AO22X1 U197 ( .IN1(n1127), .IN2(N291), .IN3(\regfile[4][1] ), .IN4(n1122), 
        .Q(n317) );
  AO22X1 U198 ( .IN1(n1126), .IN2(N309), .IN3(\regfile[4][19] ), .IN4(n1122), 
        .Q(n335) );
  AO22X1 U199 ( .IN1(n1126), .IN2(N308), .IN3(\regfile[4][18] ), .IN4(n1122), 
        .Q(n334) );
  AO22X1 U200 ( .IN1(n1126), .IN2(N307), .IN3(\regfile[4][17] ), .IN4(n1122), 
        .Q(n333) );
  AO22X1 U201 ( .IN1(n1126), .IN2(N306), .IN3(\regfile[4][16] ), .IN4(n1122), 
        .Q(n332) );
  AO22X1 U202 ( .IN1(n1126), .IN2(N305), .IN3(\regfile[4][15] ), .IN4(n1122), 
        .Q(n331) );
  AO22X1 U203 ( .IN1(n1126), .IN2(N304), .IN3(\regfile[4][14] ), .IN4(n1122), 
        .Q(n330) );
  AO22X1 U204 ( .IN1(n1126), .IN2(N303), .IN3(\regfile[4][13] ), .IN4(n1122), 
        .Q(n329) );
  AO22X1 U205 ( .IN1(n1125), .IN2(N302), .IN3(\regfile[4][12] ), .IN4(n1122), 
        .Q(n328) );
  AO22X1 U206 ( .IN1(n1125), .IN2(N301), .IN3(\regfile[4][11] ), .IN4(n1122), 
        .Q(n327) );
  AO22X1 U207 ( .IN1(n1125), .IN2(N300), .IN3(\regfile[4][10] ), .IN4(n1122), 
        .Q(n326) );
  AO22X1 U208 ( .IN1(n1125), .IN2(N290), .IN3(\regfile[4][0] ), .IN4(n1122), 
        .Q(n316) );
  AO22X1 U212 ( .IN1(n1121), .IN2(N299), .IN3(\regfile[3][9] ), .IN4(n1116), 
        .Q(n293) );
  AO22X1 U213 ( .IN1(n1121), .IN2(N298), .IN3(\regfile[3][8] ), .IN4(n1116), 
        .Q(n292) );
  AO22X1 U214 ( .IN1(n1121), .IN2(N297), .IN3(\regfile[3][7] ), .IN4(n1116), 
        .Q(n291) );
  AO22X1 U215 ( .IN1(n1121), .IN2(N296), .IN3(\regfile[3][6] ), .IN4(n1116), 
        .Q(n290) );
  AO22X1 U216 ( .IN1(n1121), .IN2(N295), .IN3(\regfile[3][5] ), .IN4(n1116), 
        .Q(n289) );
  AO22X1 U217 ( .IN1(n1121), .IN2(N294), .IN3(\regfile[3][4] ), .IN4(n1116), 
        .Q(n288) );
  AO22X1 U218 ( .IN1(n1121), .IN2(N293), .IN3(\regfile[3][3] ), .IN4(n1116), 
        .Q(n287) );
  AO22X1 U219 ( .IN1(n1120), .IN2(N321), .IN3(\regfile[3][31] ), .IN4(n1116), 
        .Q(n315) );
  AO22X1 U220 ( .IN1(n1120), .IN2(N320), .IN3(\regfile[3][30] ), .IN4(n1115), 
        .Q(n314) );
  AO22X1 U221 ( .IN1(n1120), .IN2(N292), .IN3(\regfile[3][2] ), .IN4(n1115), 
        .Q(n286) );
  AO22X1 U222 ( .IN1(n1120), .IN2(N319), .IN3(\regfile[3][29] ), .IN4(n1115), 
        .Q(n313) );
  AO22X1 U223 ( .IN1(n1120), .IN2(N318), .IN3(\regfile[3][28] ), .IN4(n1115), 
        .Q(n312) );
  AO22X1 U224 ( .IN1(n1120), .IN2(N317), .IN3(\regfile[3][27] ), .IN4(n1115), 
        .Q(n311) );
  AO22X1 U225 ( .IN1(n1120), .IN2(N316), .IN3(\regfile[3][26] ), .IN4(n1115), 
        .Q(n310) );
  AO22X1 U226 ( .IN1(n1119), .IN2(N315), .IN3(\regfile[3][25] ), .IN4(n1115), 
        .Q(n309) );
  AO22X1 U227 ( .IN1(n1119), .IN2(N314), .IN3(\regfile[3][24] ), .IN4(n1115), 
        .Q(n308) );
  AO22X1 U228 ( .IN1(n1119), .IN2(N313), .IN3(\regfile[3][23] ), .IN4(n1115), 
        .Q(n307) );
  AO22X1 U229 ( .IN1(n1119), .IN2(N312), .IN3(\regfile[3][22] ), .IN4(n1115), 
        .Q(n306) );
  AO22X1 U230 ( .IN1(n1119), .IN2(N311), .IN3(\regfile[3][21] ), .IN4(n1115), 
        .Q(n305) );
  AO22X1 U231 ( .IN1(n1119), .IN2(N310), .IN3(\regfile[3][20] ), .IN4(n1115), 
        .Q(n304) );
  AO22X1 U232 ( .IN1(n1119), .IN2(N291), .IN3(\regfile[3][1] ), .IN4(n1114), 
        .Q(n285) );
  AO22X1 U233 ( .IN1(n1118), .IN2(N309), .IN3(\regfile[3][19] ), .IN4(n1114), 
        .Q(n303) );
  AO22X1 U234 ( .IN1(n1118), .IN2(N308), .IN3(\regfile[3][18] ), .IN4(n1114), 
        .Q(n302) );
  AO22X1 U235 ( .IN1(n1118), .IN2(N307), .IN3(\regfile[3][17] ), .IN4(n1114), 
        .Q(n301) );
  AO22X1 U236 ( .IN1(n1118), .IN2(N306), .IN3(\regfile[3][16] ), .IN4(n1114), 
        .Q(n300) );
  AO22X1 U237 ( .IN1(n1118), .IN2(N305), .IN3(\regfile[3][15] ), .IN4(n1114), 
        .Q(n299) );
  AO22X1 U238 ( .IN1(n1118), .IN2(N304), .IN3(\regfile[3][14] ), .IN4(n1114), 
        .Q(n298) );
  AO22X1 U239 ( .IN1(n1118), .IN2(N303), .IN3(\regfile[3][13] ), .IN4(n1114), 
        .Q(n297) );
  AO22X1 U240 ( .IN1(n1117), .IN2(N302), .IN3(\regfile[3][12] ), .IN4(n1114), 
        .Q(n296) );
  AO22X1 U241 ( .IN1(n1117), .IN2(N301), .IN3(\regfile[3][11] ), .IN4(n1114), 
        .Q(n295) );
  AO22X1 U242 ( .IN1(n1117), .IN2(N300), .IN3(\regfile[3][10] ), .IN4(n1114), 
        .Q(n294) );
  AO22X1 U243 ( .IN1(n1117), .IN2(N290), .IN3(\regfile[3][0] ), .IN4(n1114), 
        .Q(n284) );
  AO22X1 U246 ( .IN1(n1113), .IN2(N299), .IN3(\regfile[2][9] ), .IN4(n1108), 
        .Q(n261) );
  AO22X1 U247 ( .IN1(n1113), .IN2(N298), .IN3(\regfile[2][8] ), .IN4(n1108), 
        .Q(n260) );
  AO22X1 U248 ( .IN1(n1113), .IN2(N297), .IN3(\regfile[2][7] ), .IN4(n1108), 
        .Q(n259) );
  AO22X1 U249 ( .IN1(n1113), .IN2(N296), .IN3(\regfile[2][6] ), .IN4(n1108), 
        .Q(n258) );
  AO22X1 U250 ( .IN1(n1113), .IN2(N295), .IN3(\regfile[2][5] ), .IN4(n1108), 
        .Q(n257) );
  AO22X1 U251 ( .IN1(n1113), .IN2(N294), .IN3(\regfile[2][4] ), .IN4(n1108), 
        .Q(n256) );
  AO22X1 U252 ( .IN1(n1113), .IN2(N293), .IN3(\regfile[2][3] ), .IN4(n1108), 
        .Q(n255) );
  AO22X1 U253 ( .IN1(n1112), .IN2(N321), .IN3(\regfile[2][31] ), .IN4(n1108), 
        .Q(n283) );
  AO22X1 U254 ( .IN1(n1112), .IN2(N320), .IN3(\regfile[2][30] ), .IN4(n1107), 
        .Q(n282) );
  AO22X1 U255 ( .IN1(n1112), .IN2(N292), .IN3(\regfile[2][2] ), .IN4(n1107), 
        .Q(n254) );
  AO22X1 U256 ( .IN1(n1112), .IN2(N319), .IN3(\regfile[2][29] ), .IN4(n1107), 
        .Q(n281) );
  AO22X1 U257 ( .IN1(n1112), .IN2(N318), .IN3(\regfile[2][28] ), .IN4(n1107), 
        .Q(n280) );
  AO22X1 U258 ( .IN1(n1112), .IN2(N317), .IN3(\regfile[2][27] ), .IN4(n1107), 
        .Q(n279) );
  AO22X1 U259 ( .IN1(n1112), .IN2(N316), .IN3(\regfile[2][26] ), .IN4(n1107), 
        .Q(n278) );
  AO22X1 U260 ( .IN1(n1111), .IN2(N315), .IN3(\regfile[2][25] ), .IN4(n1107), 
        .Q(n277) );
  AO22X1 U261 ( .IN1(n1111), .IN2(N314), .IN3(\regfile[2][24] ), .IN4(n1107), 
        .Q(n276) );
  AO22X1 U262 ( .IN1(n1111), .IN2(N313), .IN3(\regfile[2][23] ), .IN4(n1107), 
        .Q(n275) );
  AO22X1 U263 ( .IN1(n1111), .IN2(N312), .IN3(\regfile[2][22] ), .IN4(n1107), 
        .Q(n274) );
  AO22X1 U264 ( .IN1(n1111), .IN2(N311), .IN3(\regfile[2][21] ), .IN4(n1107), 
        .Q(n273) );
  AO22X1 U265 ( .IN1(n1111), .IN2(N310), .IN3(\regfile[2][20] ), .IN4(n1107), 
        .Q(n272) );
  AO22X1 U266 ( .IN1(n1111), .IN2(N291), .IN3(\regfile[2][1] ), .IN4(n1106), 
        .Q(n253) );
  AO22X1 U267 ( .IN1(n1110), .IN2(N309), .IN3(\regfile[2][19] ), .IN4(n1106), 
        .Q(n271) );
  AO22X1 U268 ( .IN1(n1110), .IN2(N308), .IN3(\regfile[2][18] ), .IN4(n1106), 
        .Q(n270) );
  AO22X1 U269 ( .IN1(n1110), .IN2(N307), .IN3(\regfile[2][17] ), .IN4(n1106), 
        .Q(n269) );
  AO22X1 U270 ( .IN1(n1110), .IN2(N306), .IN3(\regfile[2][16] ), .IN4(n1106), 
        .Q(n268) );
  AO22X1 U271 ( .IN1(n1110), .IN2(N305), .IN3(\regfile[2][15] ), .IN4(n1106), 
        .Q(n267) );
  AO22X1 U272 ( .IN1(n1110), .IN2(N304), .IN3(\regfile[2][14] ), .IN4(n1106), 
        .Q(n266) );
  AO22X1 U273 ( .IN1(n1110), .IN2(N303), .IN3(\regfile[2][13] ), .IN4(n1106), 
        .Q(n265) );
  AO22X1 U274 ( .IN1(n1109), .IN2(N302), .IN3(\regfile[2][12] ), .IN4(n1106), 
        .Q(n264) );
  AO22X1 U275 ( .IN1(n1109), .IN2(N301), .IN3(\regfile[2][11] ), .IN4(n1106), 
        .Q(n263) );
  AO22X1 U276 ( .IN1(n1109), .IN2(N300), .IN3(\regfile[2][10] ), .IN4(n1106), 
        .Q(n262) );
  AO22X1 U277 ( .IN1(n1109), .IN2(N290), .IN3(\regfile[2][0] ), .IN4(n1106), 
        .Q(n252) );
  AO22X1 U280 ( .IN1(n1105), .IN2(N299), .IN3(\regfile[1][9] ), .IN4(n1100), 
        .Q(n229) );
  AO22X1 U281 ( .IN1(n1105), .IN2(N298), .IN3(\regfile[1][8] ), .IN4(n1100), 
        .Q(n228) );
  AO22X1 U282 ( .IN1(n1105), .IN2(N297), .IN3(\regfile[1][7] ), .IN4(n1100), 
        .Q(n227) );
  AO22X1 U283 ( .IN1(n1105), .IN2(N296), .IN3(\regfile[1][6] ), .IN4(n1100), 
        .Q(n226) );
  AO22X1 U284 ( .IN1(n1105), .IN2(N295), .IN3(\regfile[1][5] ), .IN4(n1100), 
        .Q(n225) );
  AO22X1 U285 ( .IN1(n1105), .IN2(N294), .IN3(\regfile[1][4] ), .IN4(n1100), 
        .Q(n224) );
  AO22X1 U286 ( .IN1(n1105), .IN2(N293), .IN3(\regfile[1][3] ), .IN4(n1100), 
        .Q(n223) );
  AO22X1 U287 ( .IN1(n1104), .IN2(N321), .IN3(\regfile[1][31] ), .IN4(n1100), 
        .Q(n251) );
  AO22X1 U288 ( .IN1(n1104), .IN2(N320), .IN3(\regfile[1][30] ), .IN4(n1099), 
        .Q(n250) );
  AO22X1 U289 ( .IN1(n1104), .IN2(N292), .IN3(\regfile[1][2] ), .IN4(n1099), 
        .Q(n222) );
  AO22X1 U290 ( .IN1(n1104), .IN2(N319), .IN3(\regfile[1][29] ), .IN4(n1099), 
        .Q(n249) );
  AO22X1 U291 ( .IN1(n1104), .IN2(N318), .IN3(\regfile[1][28] ), .IN4(n1099), 
        .Q(n248) );
  AO22X1 U292 ( .IN1(n1104), .IN2(N317), .IN3(\regfile[1][27] ), .IN4(n1099), 
        .Q(n247) );
  AO22X1 U293 ( .IN1(n1104), .IN2(N316), .IN3(\regfile[1][26] ), .IN4(n1099), 
        .Q(n246) );
  AO22X1 U294 ( .IN1(n1103), .IN2(N315), .IN3(\regfile[1][25] ), .IN4(n1099), 
        .Q(n245) );
  AO22X1 U295 ( .IN1(n1103), .IN2(N314), .IN3(\regfile[1][24] ), .IN4(n1099), 
        .Q(n244) );
  AO22X1 U296 ( .IN1(n1103), .IN2(N313), .IN3(\regfile[1][23] ), .IN4(n1099), 
        .Q(n243) );
  AO22X1 U297 ( .IN1(n1103), .IN2(N312), .IN3(\regfile[1][22] ), .IN4(n1099), 
        .Q(n242) );
  AO22X1 U298 ( .IN1(n1103), .IN2(N311), .IN3(\regfile[1][21] ), .IN4(n1099), 
        .Q(n241) );
  AO22X1 U299 ( .IN1(n1103), .IN2(N310), .IN3(\regfile[1][20] ), .IN4(n1099), 
        .Q(n240) );
  AO22X1 U300 ( .IN1(n1103), .IN2(N291), .IN3(\regfile[1][1] ), .IN4(n1098), 
        .Q(n221) );
  AO22X1 U301 ( .IN1(n1102), .IN2(N309), .IN3(\regfile[1][19] ), .IN4(n1098), 
        .Q(n239) );
  AO22X1 U302 ( .IN1(n1102), .IN2(N308), .IN3(\regfile[1][18] ), .IN4(n1098), 
        .Q(n238) );
  AO22X1 U303 ( .IN1(n1102), .IN2(N307), .IN3(\regfile[1][17] ), .IN4(n1098), 
        .Q(n237) );
  AO22X1 U304 ( .IN1(n1102), .IN2(N306), .IN3(\regfile[1][16] ), .IN4(n1098), 
        .Q(n236) );
  AO22X1 U305 ( .IN1(n1102), .IN2(N305), .IN3(\regfile[1][15] ), .IN4(n1098), 
        .Q(n235) );
  AO22X1 U306 ( .IN1(n1102), .IN2(N304), .IN3(\regfile[1][14] ), .IN4(n1098), 
        .Q(n234) );
  AO22X1 U307 ( .IN1(n1102), .IN2(N303), .IN3(\regfile[1][13] ), .IN4(n1098), 
        .Q(n233) );
  AO22X1 U308 ( .IN1(n1101), .IN2(N302), .IN3(\regfile[1][12] ), .IN4(n1098), 
        .Q(n232) );
  AO22X1 U309 ( .IN1(n1101), .IN2(N301), .IN3(\regfile[1][11] ), .IN4(n1098), 
        .Q(n231) );
  AO22X1 U310 ( .IN1(n1101), .IN2(N300), .IN3(\regfile[1][10] ), .IN4(n1098), 
        .Q(n230) );
  AO22X1 U311 ( .IN1(n1101), .IN2(N290), .IN3(\regfile[1][0] ), .IN4(n1098), 
        .Q(n220) );
  AO22X1 U314 ( .IN1(n1097), .IN2(N299), .IN3(\regfile[15][9] ), .IN4(n1092), 
        .Q(n677) );
  AO22X1 U315 ( .IN1(n1097), .IN2(N298), .IN3(\regfile[15][8] ), .IN4(n1092), 
        .Q(n676) );
  AO22X1 U316 ( .IN1(n1097), .IN2(N297), .IN3(\regfile[15][7] ), .IN4(n1092), 
        .Q(n675) );
  AO22X1 U317 ( .IN1(n1097), .IN2(N296), .IN3(\regfile[15][6] ), .IN4(n1092), 
        .Q(n674) );
  AO22X1 U318 ( .IN1(n1097), .IN2(N295), .IN3(\regfile[15][5] ), .IN4(n1092), 
        .Q(n673) );
  AO22X1 U319 ( .IN1(n1097), .IN2(N294), .IN3(\regfile[15][4] ), .IN4(n1092), 
        .Q(n672) );
  AO22X1 U320 ( .IN1(n1097), .IN2(N293), .IN3(\regfile[15][3] ), .IN4(n1092), 
        .Q(n671) );
  AO22X1 U321 ( .IN1(n1096), .IN2(N321), .IN3(\regfile[15][31] ), .IN4(n1092), 
        .Q(n699) );
  AO22X1 U322 ( .IN1(n1096), .IN2(N320), .IN3(\regfile[15][30] ), .IN4(n1091), 
        .Q(n698) );
  AO22X1 U323 ( .IN1(n1096), .IN2(N292), .IN3(\regfile[15][2] ), .IN4(n1091), 
        .Q(n670) );
  AO22X1 U324 ( .IN1(n1096), .IN2(N319), .IN3(\regfile[15][29] ), .IN4(n1091), 
        .Q(n697) );
  AO22X1 U325 ( .IN1(n1096), .IN2(N318), .IN3(\regfile[15][28] ), .IN4(n1091), 
        .Q(n696) );
  AO22X1 U326 ( .IN1(n1096), .IN2(N317), .IN3(\regfile[15][27] ), .IN4(n1091), 
        .Q(n695) );
  AO22X1 U327 ( .IN1(n1096), .IN2(N316), .IN3(\regfile[15][26] ), .IN4(n1091), 
        .Q(n694) );
  AO22X1 U328 ( .IN1(n1095), .IN2(N315), .IN3(\regfile[15][25] ), .IN4(n1091), 
        .Q(n693) );
  AO22X1 U329 ( .IN1(n1095), .IN2(N314), .IN3(\regfile[15][24] ), .IN4(n1091), 
        .Q(n692) );
  AO22X1 U330 ( .IN1(n1095), .IN2(N313), .IN3(\regfile[15][23] ), .IN4(n1091), 
        .Q(n691) );
  AO22X1 U331 ( .IN1(n1095), .IN2(N312), .IN3(\regfile[15][22] ), .IN4(n1091), 
        .Q(n690) );
  AO22X1 U332 ( .IN1(n1095), .IN2(N311), .IN3(\regfile[15][21] ), .IN4(n1091), 
        .Q(n689) );
  AO22X1 U333 ( .IN1(n1095), .IN2(N310), .IN3(\regfile[15][20] ), .IN4(n1091), 
        .Q(n688) );
  AO22X1 U334 ( .IN1(n1095), .IN2(N291), .IN3(\regfile[15][1] ), .IN4(n1090), 
        .Q(n669) );
  AO22X1 U335 ( .IN1(n1094), .IN2(N309), .IN3(\regfile[15][19] ), .IN4(n1090), 
        .Q(n687) );
  AO22X1 U336 ( .IN1(n1094), .IN2(N308), .IN3(\regfile[15][18] ), .IN4(n1090), 
        .Q(n686) );
  AO22X1 U337 ( .IN1(n1094), .IN2(N307), .IN3(\regfile[15][17] ), .IN4(n1090), 
        .Q(n685) );
  AO22X1 U338 ( .IN1(n1094), .IN2(N306), .IN3(\regfile[15][16] ), .IN4(n1090), 
        .Q(n684) );
  AO22X1 U339 ( .IN1(n1094), .IN2(N305), .IN3(\regfile[15][15] ), .IN4(n1090), 
        .Q(n683) );
  AO22X1 U340 ( .IN1(n1094), .IN2(N304), .IN3(\regfile[15][14] ), .IN4(n1090), 
        .Q(n682) );
  AO22X1 U341 ( .IN1(n1094), .IN2(N303), .IN3(\regfile[15][13] ), .IN4(n1090), 
        .Q(n681) );
  AO22X1 U342 ( .IN1(n1093), .IN2(N302), .IN3(\regfile[15][12] ), .IN4(n1090), 
        .Q(n680) );
  AO22X1 U343 ( .IN1(n1093), .IN2(N301), .IN3(\regfile[15][11] ), .IN4(n1090), 
        .Q(n679) );
  AO22X1 U344 ( .IN1(n1093), .IN2(N300), .IN3(\regfile[15][10] ), .IN4(n1090), 
        .Q(n678) );
  AO22X1 U345 ( .IN1(n1093), .IN2(N290), .IN3(\regfile[15][0] ), .IN4(n1090), 
        .Q(n668) );
  AO22X1 U348 ( .IN1(n1089), .IN2(N299), .IN3(\regfile[14][9] ), .IN4(n1084), 
        .Q(n645) );
  AO22X1 U349 ( .IN1(n1089), .IN2(N298), .IN3(\regfile[14][8] ), .IN4(n1084), 
        .Q(n644) );
  AO22X1 U350 ( .IN1(n1089), .IN2(N297), .IN3(\regfile[14][7] ), .IN4(n1084), 
        .Q(n643) );
  AO22X1 U351 ( .IN1(n1089), .IN2(N296), .IN3(\regfile[14][6] ), .IN4(n1084), 
        .Q(n642) );
  AO22X1 U352 ( .IN1(n1089), .IN2(N295), .IN3(\regfile[14][5] ), .IN4(n1084), 
        .Q(n641) );
  AO22X1 U353 ( .IN1(n1089), .IN2(N294), .IN3(\regfile[14][4] ), .IN4(n1084), 
        .Q(n640) );
  AO22X1 U354 ( .IN1(n1089), .IN2(N293), .IN3(\regfile[14][3] ), .IN4(n1084), 
        .Q(n639) );
  AO22X1 U355 ( .IN1(n1088), .IN2(N321), .IN3(\regfile[14][31] ), .IN4(n1084), 
        .Q(n667) );
  AO22X1 U356 ( .IN1(n1088), .IN2(N320), .IN3(\regfile[14][30] ), .IN4(n1083), 
        .Q(n666) );
  AO22X1 U357 ( .IN1(n1088), .IN2(N292), .IN3(\regfile[14][2] ), .IN4(n1083), 
        .Q(n638) );
  AO22X1 U358 ( .IN1(n1088), .IN2(N319), .IN3(\regfile[14][29] ), .IN4(n1083), 
        .Q(n665) );
  AO22X1 U359 ( .IN1(n1088), .IN2(N318), .IN3(\regfile[14][28] ), .IN4(n1083), 
        .Q(n664) );
  AO22X1 U360 ( .IN1(n1088), .IN2(N317), .IN3(\regfile[14][27] ), .IN4(n1083), 
        .Q(n663) );
  AO22X1 U361 ( .IN1(n1088), .IN2(N316), .IN3(\regfile[14][26] ), .IN4(n1083), 
        .Q(n662) );
  AO22X1 U362 ( .IN1(n1087), .IN2(N315), .IN3(\regfile[14][25] ), .IN4(n1083), 
        .Q(n661) );
  AO22X1 U363 ( .IN1(n1087), .IN2(N314), .IN3(\regfile[14][24] ), .IN4(n1083), 
        .Q(n660) );
  AO22X1 U364 ( .IN1(n1087), .IN2(N313), .IN3(\regfile[14][23] ), .IN4(n1083), 
        .Q(n659) );
  AO22X1 U365 ( .IN1(n1087), .IN2(N312), .IN3(\regfile[14][22] ), .IN4(n1083), 
        .Q(n658) );
  AO22X1 U366 ( .IN1(n1087), .IN2(N311), .IN3(\regfile[14][21] ), .IN4(n1083), 
        .Q(n657) );
  AO22X1 U367 ( .IN1(n1087), .IN2(N310), .IN3(\regfile[14][20] ), .IN4(n1083), 
        .Q(n656) );
  AO22X1 U368 ( .IN1(n1087), .IN2(N291), .IN3(\regfile[14][1] ), .IN4(n1082), 
        .Q(n637) );
  AO22X1 U369 ( .IN1(n1086), .IN2(N309), .IN3(\regfile[14][19] ), .IN4(n1082), 
        .Q(n655) );
  AO22X1 U370 ( .IN1(n1086), .IN2(N308), .IN3(\regfile[14][18] ), .IN4(n1082), 
        .Q(n654) );
  AO22X1 U371 ( .IN1(n1086), .IN2(N307), .IN3(\regfile[14][17] ), .IN4(n1082), 
        .Q(n653) );
  AO22X1 U372 ( .IN1(n1086), .IN2(N306), .IN3(\regfile[14][16] ), .IN4(n1082), 
        .Q(n652) );
  AO22X1 U373 ( .IN1(n1086), .IN2(N305), .IN3(\regfile[14][15] ), .IN4(n1082), 
        .Q(n651) );
  AO22X1 U374 ( .IN1(n1086), .IN2(N304), .IN3(\regfile[14][14] ), .IN4(n1082), 
        .Q(n650) );
  AO22X1 U375 ( .IN1(n1086), .IN2(N303), .IN3(\regfile[14][13] ), .IN4(n1082), 
        .Q(n649) );
  AO22X1 U376 ( .IN1(n1085), .IN2(N302), .IN3(\regfile[14][12] ), .IN4(n1082), 
        .Q(n648) );
  AO22X1 U377 ( .IN1(n1085), .IN2(N301), .IN3(\regfile[14][11] ), .IN4(n1082), 
        .Q(n647) );
  AO22X1 U378 ( .IN1(n1085), .IN2(N300), .IN3(\regfile[14][10] ), .IN4(n1082), 
        .Q(n646) );
  AO22X1 U379 ( .IN1(n1085), .IN2(N290), .IN3(\regfile[14][0] ), .IN4(n1082), 
        .Q(n636) );
  AO22X1 U382 ( .IN1(n1081), .IN2(N299), .IN3(\regfile[13][9] ), .IN4(n1076), 
        .Q(n613) );
  AO22X1 U383 ( .IN1(n1081), .IN2(N298), .IN3(\regfile[13][8] ), .IN4(n1076), 
        .Q(n612) );
  AO22X1 U384 ( .IN1(n1081), .IN2(N297), .IN3(\regfile[13][7] ), .IN4(n1076), 
        .Q(n611) );
  AO22X1 U385 ( .IN1(n1081), .IN2(N296), .IN3(\regfile[13][6] ), .IN4(n1076), 
        .Q(n610) );
  AO22X1 U386 ( .IN1(n1081), .IN2(N295), .IN3(\regfile[13][5] ), .IN4(n1076), 
        .Q(n609) );
  AO22X1 U387 ( .IN1(n1081), .IN2(N294), .IN3(\regfile[13][4] ), .IN4(n1076), 
        .Q(n608) );
  AO22X1 U388 ( .IN1(n1081), .IN2(N293), .IN3(\regfile[13][3] ), .IN4(n1076), 
        .Q(n607) );
  AO22X1 U389 ( .IN1(n1080), .IN2(N321), .IN3(\regfile[13][31] ), .IN4(n1076), 
        .Q(n635) );
  AO22X1 U390 ( .IN1(n1080), .IN2(N320), .IN3(\regfile[13][30] ), .IN4(n1075), 
        .Q(n634) );
  AO22X1 U391 ( .IN1(n1080), .IN2(N292), .IN3(\regfile[13][2] ), .IN4(n1075), 
        .Q(n606) );
  AO22X1 U392 ( .IN1(n1080), .IN2(N319), .IN3(\regfile[13][29] ), .IN4(n1075), 
        .Q(n633) );
  AO22X1 U393 ( .IN1(n1080), .IN2(N318), .IN3(\regfile[13][28] ), .IN4(n1075), 
        .Q(n632) );
  AO22X1 U394 ( .IN1(n1080), .IN2(N317), .IN3(\regfile[13][27] ), .IN4(n1075), 
        .Q(n631) );
  AO22X1 U395 ( .IN1(n1080), .IN2(N316), .IN3(\regfile[13][26] ), .IN4(n1075), 
        .Q(n630) );
  AO22X1 U396 ( .IN1(n1079), .IN2(N315), .IN3(\regfile[13][25] ), .IN4(n1075), 
        .Q(n629) );
  AO22X1 U397 ( .IN1(n1079), .IN2(N314), .IN3(\regfile[13][24] ), .IN4(n1075), 
        .Q(n628) );
  AO22X1 U398 ( .IN1(n1079), .IN2(N313), .IN3(\regfile[13][23] ), .IN4(n1075), 
        .Q(n627) );
  AO22X1 U399 ( .IN1(n1079), .IN2(N312), .IN3(\regfile[13][22] ), .IN4(n1075), 
        .Q(n626) );
  AO22X1 U400 ( .IN1(n1079), .IN2(N311), .IN3(\regfile[13][21] ), .IN4(n1075), 
        .Q(n625) );
  AO22X1 U401 ( .IN1(n1079), .IN2(N310), .IN3(\regfile[13][20] ), .IN4(n1075), 
        .Q(n624) );
  AO22X1 U402 ( .IN1(n1079), .IN2(N291), .IN3(\regfile[13][1] ), .IN4(n1074), 
        .Q(n605) );
  AO22X1 U403 ( .IN1(n1078), .IN2(N309), .IN3(\regfile[13][19] ), .IN4(n1074), 
        .Q(n623) );
  AO22X1 U404 ( .IN1(n1078), .IN2(N308), .IN3(\regfile[13][18] ), .IN4(n1074), 
        .Q(n622) );
  AO22X1 U405 ( .IN1(n1078), .IN2(N307), .IN3(\regfile[13][17] ), .IN4(n1074), 
        .Q(n621) );
  AO22X1 U406 ( .IN1(n1078), .IN2(N306), .IN3(\regfile[13][16] ), .IN4(n1074), 
        .Q(n620) );
  AO22X1 U407 ( .IN1(n1078), .IN2(N305), .IN3(\regfile[13][15] ), .IN4(n1074), 
        .Q(n619) );
  AO22X1 U408 ( .IN1(n1078), .IN2(N304), .IN3(\regfile[13][14] ), .IN4(n1074), 
        .Q(n618) );
  AO22X1 U409 ( .IN1(n1078), .IN2(N303), .IN3(\regfile[13][13] ), .IN4(n1074), 
        .Q(n617) );
  AO22X1 U410 ( .IN1(n1077), .IN2(N302), .IN3(\regfile[13][12] ), .IN4(n1074), 
        .Q(n616) );
  AO22X1 U411 ( .IN1(n1077), .IN2(N301), .IN3(\regfile[13][11] ), .IN4(n1074), 
        .Q(n615) );
  AO22X1 U412 ( .IN1(n1077), .IN2(N300), .IN3(\regfile[13][10] ), .IN4(n1074), 
        .Q(n614) );
  AO22X1 U413 ( .IN1(n1077), .IN2(N290), .IN3(\regfile[13][0] ), .IN4(n1074), 
        .Q(n604) );
  AO22X1 U417 ( .IN1(n1073), .IN2(N299), .IN3(\regfile[12][9] ), .IN4(n1068), 
        .Q(n581) );
  AO22X1 U418 ( .IN1(n1073), .IN2(N298), .IN3(\regfile[12][8] ), .IN4(n1068), 
        .Q(n580) );
  AO22X1 U419 ( .IN1(n1073), .IN2(N297), .IN3(\regfile[12][7] ), .IN4(n1068), 
        .Q(n579) );
  AO22X1 U420 ( .IN1(n1073), .IN2(N296), .IN3(\regfile[12][6] ), .IN4(n1068), 
        .Q(n578) );
  AO22X1 U421 ( .IN1(n1073), .IN2(N295), .IN3(\regfile[12][5] ), .IN4(n1068), 
        .Q(n577) );
  AO22X1 U422 ( .IN1(n1073), .IN2(N294), .IN3(\regfile[12][4] ), .IN4(n1068), 
        .Q(n576) );
  AO22X1 U423 ( .IN1(n1073), .IN2(N293), .IN3(\regfile[12][3] ), .IN4(n1068), 
        .Q(n575) );
  AO22X1 U424 ( .IN1(n1072), .IN2(N321), .IN3(\regfile[12][31] ), .IN4(n1068), 
        .Q(n603) );
  AO22X1 U425 ( .IN1(n1072), .IN2(N320), .IN3(\regfile[12][30] ), .IN4(n1067), 
        .Q(n602) );
  AO22X1 U426 ( .IN1(n1072), .IN2(N292), .IN3(\regfile[12][2] ), .IN4(n1067), 
        .Q(n574) );
  AO22X1 U427 ( .IN1(n1072), .IN2(N319), .IN3(\regfile[12][29] ), .IN4(n1067), 
        .Q(n601) );
  AO22X1 U428 ( .IN1(n1072), .IN2(N318), .IN3(\regfile[12][28] ), .IN4(n1067), 
        .Q(n600) );
  AO22X1 U429 ( .IN1(n1072), .IN2(N317), .IN3(\regfile[12][27] ), .IN4(n1067), 
        .Q(n599) );
  AO22X1 U430 ( .IN1(n1072), .IN2(N316), .IN3(\regfile[12][26] ), .IN4(n1067), 
        .Q(n598) );
  AO22X1 U431 ( .IN1(n1071), .IN2(N315), .IN3(\regfile[12][25] ), .IN4(n1067), 
        .Q(n597) );
  AO22X1 U432 ( .IN1(n1071), .IN2(N314), .IN3(\regfile[12][24] ), .IN4(n1067), 
        .Q(n596) );
  AO22X1 U433 ( .IN1(n1071), .IN2(N313), .IN3(\regfile[12][23] ), .IN4(n1067), 
        .Q(n595) );
  AO22X1 U434 ( .IN1(n1071), .IN2(N312), .IN3(\regfile[12][22] ), .IN4(n1067), 
        .Q(n594) );
  AO22X1 U435 ( .IN1(n1071), .IN2(N311), .IN3(\regfile[12][21] ), .IN4(n1067), 
        .Q(n593) );
  AO22X1 U436 ( .IN1(n1071), .IN2(N310), .IN3(\regfile[12][20] ), .IN4(n1067), 
        .Q(n592) );
  AO22X1 U437 ( .IN1(n1071), .IN2(N291), .IN3(\regfile[12][1] ), .IN4(n1066), 
        .Q(n573) );
  AO22X1 U438 ( .IN1(n1070), .IN2(N309), .IN3(\regfile[12][19] ), .IN4(n1066), 
        .Q(n591) );
  AO22X1 U439 ( .IN1(n1070), .IN2(N308), .IN3(\regfile[12][18] ), .IN4(n1066), 
        .Q(n590) );
  AO22X1 U440 ( .IN1(n1070), .IN2(N307), .IN3(\regfile[12][17] ), .IN4(n1066), 
        .Q(n589) );
  AO22X1 U441 ( .IN1(n1070), .IN2(N306), .IN3(\regfile[12][16] ), .IN4(n1066), 
        .Q(n588) );
  AO22X1 U442 ( .IN1(n1070), .IN2(N305), .IN3(\regfile[12][15] ), .IN4(n1066), 
        .Q(n587) );
  AO22X1 U443 ( .IN1(n1070), .IN2(N304), .IN3(\regfile[12][14] ), .IN4(n1066), 
        .Q(n586) );
  AO22X1 U444 ( .IN1(n1070), .IN2(N303), .IN3(\regfile[12][13] ), .IN4(n1066), 
        .Q(n585) );
  AO22X1 U445 ( .IN1(n1069), .IN2(N302), .IN3(\regfile[12][12] ), .IN4(n1066), 
        .Q(n584) );
  AO22X1 U446 ( .IN1(n1069), .IN2(N301), .IN3(\regfile[12][11] ), .IN4(n1066), 
        .Q(n583) );
  AO22X1 U447 ( .IN1(n1069), .IN2(N300), .IN3(\regfile[12][10] ), .IN4(n1066), 
        .Q(n582) );
  AO22X1 U448 ( .IN1(n1069), .IN2(N290), .IN3(\regfile[12][0] ), .IN4(n1066), 
        .Q(n572) );
  AO22X1 U452 ( .IN1(n1065), .IN2(N299), .IN3(\regfile[11][9] ), .IN4(n1060), 
        .Q(n549) );
  AO22X1 U453 ( .IN1(n1065), .IN2(N298), .IN3(\regfile[11][8] ), .IN4(n1060), 
        .Q(n548) );
  AO22X1 U454 ( .IN1(n1065), .IN2(N297), .IN3(\regfile[11][7] ), .IN4(n1060), 
        .Q(n547) );
  AO22X1 U455 ( .IN1(n1065), .IN2(N296), .IN3(\regfile[11][6] ), .IN4(n1060), 
        .Q(n546) );
  AO22X1 U456 ( .IN1(n1065), .IN2(N295), .IN3(\regfile[11][5] ), .IN4(n1060), 
        .Q(n545) );
  AO22X1 U457 ( .IN1(n1065), .IN2(N294), .IN3(\regfile[11][4] ), .IN4(n1060), 
        .Q(n544) );
  AO22X1 U458 ( .IN1(n1065), .IN2(N293), .IN3(\regfile[11][3] ), .IN4(n1060), 
        .Q(n543) );
  AO22X1 U459 ( .IN1(n1064), .IN2(N321), .IN3(\regfile[11][31] ), .IN4(n1060), 
        .Q(n571) );
  AO22X1 U460 ( .IN1(n1064), .IN2(N320), .IN3(\regfile[11][30] ), .IN4(n1059), 
        .Q(n570) );
  AO22X1 U461 ( .IN1(n1064), .IN2(N292), .IN3(\regfile[11][2] ), .IN4(n1059), 
        .Q(n542) );
  AO22X1 U462 ( .IN1(n1064), .IN2(N319), .IN3(\regfile[11][29] ), .IN4(n1059), 
        .Q(n569) );
  AO22X1 U463 ( .IN1(n1064), .IN2(N318), .IN3(\regfile[11][28] ), .IN4(n1059), 
        .Q(n568) );
  AO22X1 U464 ( .IN1(n1064), .IN2(N317), .IN3(\regfile[11][27] ), .IN4(n1059), 
        .Q(n567) );
  AO22X1 U465 ( .IN1(n1064), .IN2(N316), .IN3(\regfile[11][26] ), .IN4(n1059), 
        .Q(n566) );
  AO22X1 U466 ( .IN1(n1063), .IN2(N315), .IN3(\regfile[11][25] ), .IN4(n1059), 
        .Q(n565) );
  AO22X1 U467 ( .IN1(n1063), .IN2(N314), .IN3(\regfile[11][24] ), .IN4(n1059), 
        .Q(n564) );
  AO22X1 U468 ( .IN1(n1063), .IN2(N313), .IN3(\regfile[11][23] ), .IN4(n1059), 
        .Q(n563) );
  AO22X1 U469 ( .IN1(n1063), .IN2(N312), .IN3(\regfile[11][22] ), .IN4(n1059), 
        .Q(n562) );
  AO22X1 U470 ( .IN1(n1063), .IN2(N311), .IN3(\regfile[11][21] ), .IN4(n1059), 
        .Q(n561) );
  AO22X1 U471 ( .IN1(n1063), .IN2(N310), .IN3(\regfile[11][20] ), .IN4(n1059), 
        .Q(n560) );
  AO22X1 U472 ( .IN1(n1063), .IN2(N291), .IN3(\regfile[11][1] ), .IN4(n1058), 
        .Q(n541) );
  AO22X1 U473 ( .IN1(n1062), .IN2(N309), .IN3(\regfile[11][19] ), .IN4(n1058), 
        .Q(n559) );
  AO22X1 U474 ( .IN1(n1062), .IN2(N308), .IN3(\regfile[11][18] ), .IN4(n1058), 
        .Q(n558) );
  AO22X1 U475 ( .IN1(n1062), .IN2(N307), .IN3(\regfile[11][17] ), .IN4(n1058), 
        .Q(n557) );
  AO22X1 U476 ( .IN1(n1062), .IN2(N306), .IN3(\regfile[11][16] ), .IN4(n1058), 
        .Q(n556) );
  AO22X1 U477 ( .IN1(n1062), .IN2(N305), .IN3(\regfile[11][15] ), .IN4(n1058), 
        .Q(n555) );
  AO22X1 U478 ( .IN1(n1062), .IN2(N304), .IN3(\regfile[11][14] ), .IN4(n1058), 
        .Q(n554) );
  AO22X1 U479 ( .IN1(n1062), .IN2(N303), .IN3(\regfile[11][13] ), .IN4(n1058), 
        .Q(n553) );
  AO22X1 U480 ( .IN1(n1061), .IN2(N302), .IN3(\regfile[11][12] ), .IN4(n1058), 
        .Q(n552) );
  AO22X1 U481 ( .IN1(n1061), .IN2(N301), .IN3(\regfile[11][11] ), .IN4(n1058), 
        .Q(n551) );
  AO22X1 U482 ( .IN1(n1061), .IN2(N300), .IN3(\regfile[11][10] ), .IN4(n1058), 
        .Q(n550) );
  AO22X1 U483 ( .IN1(n1061), .IN2(N290), .IN3(\regfile[11][0] ), .IN4(n1058), 
        .Q(n540) );
  AO22X1 U487 ( .IN1(n1057), .IN2(N299), .IN3(\regfile[10][9] ), .IN4(n1052), 
        .Q(n517) );
  AO22X1 U488 ( .IN1(n1057), .IN2(N298), .IN3(\regfile[10][8] ), .IN4(n1052), 
        .Q(n516) );
  AO22X1 U489 ( .IN1(n1057), .IN2(N297), .IN3(\regfile[10][7] ), .IN4(n1052), 
        .Q(n515) );
  AO22X1 U490 ( .IN1(n1057), .IN2(N296), .IN3(\regfile[10][6] ), .IN4(n1052), 
        .Q(n514) );
  AO22X1 U491 ( .IN1(n1057), .IN2(N295), .IN3(\regfile[10][5] ), .IN4(n1052), 
        .Q(n513) );
  AO22X1 U492 ( .IN1(n1057), .IN2(N294), .IN3(\regfile[10][4] ), .IN4(n1052), 
        .Q(n512) );
  AO22X1 U493 ( .IN1(n1057), .IN2(N293), .IN3(\regfile[10][3] ), .IN4(n1052), 
        .Q(n511) );
  AO22X1 U494 ( .IN1(n1056), .IN2(N321), .IN3(\regfile[10][31] ), .IN4(n1052), 
        .Q(n539) );
  AO22X1 U495 ( .IN1(n1056), .IN2(N320), .IN3(\regfile[10][30] ), .IN4(n1051), 
        .Q(n538) );
  AO22X1 U496 ( .IN1(n1056), .IN2(N292), .IN3(\regfile[10][2] ), .IN4(n1051), 
        .Q(n510) );
  AO22X1 U497 ( .IN1(n1056), .IN2(N319), .IN3(\regfile[10][29] ), .IN4(n1051), 
        .Q(n537) );
  AO22X1 U498 ( .IN1(n1056), .IN2(N318), .IN3(\regfile[10][28] ), .IN4(n1051), 
        .Q(n536) );
  AO22X1 U499 ( .IN1(n1056), .IN2(N317), .IN3(\regfile[10][27] ), .IN4(n1051), 
        .Q(n535) );
  AO22X1 U500 ( .IN1(n1056), .IN2(N316), .IN3(\regfile[10][26] ), .IN4(n1051), 
        .Q(n534) );
  AO22X1 U501 ( .IN1(n1055), .IN2(N315), .IN3(\regfile[10][25] ), .IN4(n1051), 
        .Q(n533) );
  AO22X1 U502 ( .IN1(n1055), .IN2(N314), .IN3(\regfile[10][24] ), .IN4(n1051), 
        .Q(n532) );
  AO22X1 U503 ( .IN1(n1055), .IN2(N313), .IN3(\regfile[10][23] ), .IN4(n1051), 
        .Q(n531) );
  AO22X1 U504 ( .IN1(n1055), .IN2(N312), .IN3(\regfile[10][22] ), .IN4(n1051), 
        .Q(n530) );
  AO22X1 U505 ( .IN1(n1055), .IN2(N311), .IN3(\regfile[10][21] ), .IN4(n1051), 
        .Q(n529) );
  AO22X1 U506 ( .IN1(n1055), .IN2(N310), .IN3(\regfile[10][20] ), .IN4(n1051), 
        .Q(n528) );
  AO22X1 U507 ( .IN1(n1055), .IN2(N291), .IN3(\regfile[10][1] ), .IN4(n1050), 
        .Q(n509) );
  AO22X1 U508 ( .IN1(n1054), .IN2(N309), .IN3(\regfile[10][19] ), .IN4(n1050), 
        .Q(n527) );
  AO22X1 U509 ( .IN1(n1054), .IN2(N308), .IN3(\regfile[10][18] ), .IN4(n1050), 
        .Q(n526) );
  AO22X1 U510 ( .IN1(n1054), .IN2(N307), .IN3(\regfile[10][17] ), .IN4(n1050), 
        .Q(n525) );
  AO22X1 U511 ( .IN1(n1054), .IN2(N306), .IN3(\regfile[10][16] ), .IN4(n1050), 
        .Q(n524) );
  AO22X1 U512 ( .IN1(n1054), .IN2(N305), .IN3(\regfile[10][15] ), .IN4(n1050), 
        .Q(n523) );
  AO22X1 U513 ( .IN1(n1054), .IN2(N304), .IN3(\regfile[10][14] ), .IN4(n1050), 
        .Q(n522) );
  AO22X1 U514 ( .IN1(n1054), .IN2(N303), .IN3(\regfile[10][13] ), .IN4(n1050), 
        .Q(n521) );
  AO22X1 U515 ( .IN1(n1053), .IN2(N302), .IN3(\regfile[10][12] ), .IN4(n1050), 
        .Q(n520) );
  AO22X1 U516 ( .IN1(n1053), .IN2(N301), .IN3(\regfile[10][11] ), .IN4(n1050), 
        .Q(n519) );
  AO22X1 U517 ( .IN1(n1053), .IN2(N300), .IN3(\regfile[10][10] ), .IN4(n1050), 
        .Q(n518) );
  AO22X1 U518 ( .IN1(n1053), .IN2(N290), .IN3(\regfile[10][0] ), .IN4(n1050), 
        .Q(n508) );
  AO22X1 U523 ( .IN1(n1049), .IN2(N299), .IN3(\regfile[0][9] ), .IN4(n1044), 
        .Q(n197) );
  AO22X1 U524 ( .IN1(n1049), .IN2(N298), .IN3(\regfile[0][8] ), .IN4(n1044), 
        .Q(n196) );
  AO22X1 U525 ( .IN1(n1049), .IN2(N297), .IN3(\regfile[0][7] ), .IN4(n1044), 
        .Q(n195) );
  AO22X1 U526 ( .IN1(n1049), .IN2(N296), .IN3(\regfile[0][6] ), .IN4(n1044), 
        .Q(n194) );
  AO22X1 U527 ( .IN1(n1049), .IN2(N295), .IN3(\regfile[0][5] ), .IN4(n1044), 
        .Q(n193) );
  AO22X1 U528 ( .IN1(n1049), .IN2(N294), .IN3(\regfile[0][4] ), .IN4(n1044), 
        .Q(n192) );
  AO22X1 U529 ( .IN1(n1049), .IN2(N293), .IN3(\regfile[0][3] ), .IN4(n1044), 
        .Q(n191) );
  AO22X1 U530 ( .IN1(n1048), .IN2(N321), .IN3(\regfile[0][31] ), .IN4(n1044), 
        .Q(n219) );
  AO22X1 U531 ( .IN1(n1048), .IN2(N320), .IN3(\regfile[0][30] ), .IN4(n1043), 
        .Q(n218) );
  AO22X1 U532 ( .IN1(n1048), .IN2(N292), .IN3(\regfile[0][2] ), .IN4(n1043), 
        .Q(n190) );
  AO22X1 U533 ( .IN1(n1048), .IN2(N319), .IN3(\regfile[0][29] ), .IN4(n1043), 
        .Q(n217) );
  AO22X1 U534 ( .IN1(n1048), .IN2(N318), .IN3(\regfile[0][28] ), .IN4(n1043), 
        .Q(n216) );
  AO22X1 U535 ( .IN1(n1048), .IN2(N317), .IN3(\regfile[0][27] ), .IN4(n1043), 
        .Q(n215) );
  AO22X1 U536 ( .IN1(n1048), .IN2(N316), .IN3(\regfile[0][26] ), .IN4(n1043), 
        .Q(n214) );
  AO22X1 U537 ( .IN1(n1047), .IN2(N315), .IN3(\regfile[0][25] ), .IN4(n1043), 
        .Q(n213) );
  AO22X1 U538 ( .IN1(n1047), .IN2(N314), .IN3(\regfile[0][24] ), .IN4(n1043), 
        .Q(n212) );
  AO22X1 U539 ( .IN1(n1047), .IN2(N313), .IN3(\regfile[0][23] ), .IN4(n1043), 
        .Q(n211) );
  AO22X1 U540 ( .IN1(n1047), .IN2(N312), .IN3(\regfile[0][22] ), .IN4(n1043), 
        .Q(n210) );
  AO22X1 U541 ( .IN1(n1047), .IN2(N311), .IN3(\regfile[0][21] ), .IN4(n1043), 
        .Q(n209) );
  AO22X1 U542 ( .IN1(n1047), .IN2(N310), .IN3(\regfile[0][20] ), .IN4(n1043), 
        .Q(n208) );
  AO22X1 U543 ( .IN1(n1047), .IN2(N291), .IN3(\regfile[0][1] ), .IN4(n1042), 
        .Q(n189) );
  AO22X1 U544 ( .IN1(n1046), .IN2(N309), .IN3(\regfile[0][19] ), .IN4(n1042), 
        .Q(n207) );
  AO22X1 U545 ( .IN1(n1046), .IN2(N308), .IN3(\regfile[0][18] ), .IN4(n1042), 
        .Q(n206) );
  AO22X1 U546 ( .IN1(n1046), .IN2(N307), .IN3(\regfile[0][17] ), .IN4(n1042), 
        .Q(n205) );
  AO22X1 U547 ( .IN1(n1046), .IN2(N306), .IN3(\regfile[0][16] ), .IN4(n1042), 
        .Q(n204) );
  AO22X1 U548 ( .IN1(n1046), .IN2(N305), .IN3(\regfile[0][15] ), .IN4(n1042), 
        .Q(n203) );
  AO22X1 U549 ( .IN1(n1046), .IN2(N304), .IN3(\regfile[0][14] ), .IN4(n1042), 
        .Q(n202) );
  AO22X1 U550 ( .IN1(n1046), .IN2(N303), .IN3(\regfile[0][13] ), .IN4(n1042), 
        .Q(n201) );
  AO22X1 U551 ( .IN1(n1045), .IN2(N302), .IN3(\regfile[0][12] ), .IN4(n1042), 
        .Q(n200) );
  AO22X1 U552 ( .IN1(n1045), .IN2(N301), .IN3(\regfile[0][11] ), .IN4(n1042), 
        .Q(n199) );
  AO22X1 U553 ( .IN1(n1045), .IN2(N300), .IN3(\regfile[0][10] ), .IN4(n1042), 
        .Q(n198) );
  AO22X1 U554 ( .IN1(n1045), .IN2(N290), .IN3(\regfile[0][0] ), .IN4(n1042), 
        .Q(n188) );
  AND2X1 U563 ( .IN1(n53), .IN2(n54), .Q(n701) );
  NOR4X0 U564 ( .IN1(n55), .IN2(n56), .IN3(n57), .IN4(n58), .QN(n54) );
  OR4X1 U565 ( .IN1(N306), .IN2(N307), .IN3(N308), .IN4(N309), .Q(n58) );
  OR4X1 U566 ( .IN1(N310), .IN2(N311), .IN3(N312), .IN4(N313), .Q(n57) );
  OR4X1 U567 ( .IN1(N314), .IN2(N315), .IN3(N316), .IN4(N317), .Q(n56) );
  OR4X1 U568 ( .IN1(N318), .IN2(N319), .IN3(N320), .IN4(N321), .Q(n55) );
  NOR4X0 U569 ( .IN1(n59), .IN2(n60), .IN3(n61), .IN4(n62), .QN(n53) );
  OR4X1 U570 ( .IN1(N290), .IN2(N291), .IN3(N292), .IN4(N293), .Q(n62) );
  OR4X1 U571 ( .IN1(N294), .IN2(N295), .IN3(N296), .IN4(N297), .Q(n61) );
  OR4X1 U572 ( .IN1(N298), .IN2(N299), .IN3(N300), .IN4(N301), .Q(n60) );
  OR4X1 U573 ( .IN1(N302), .IN2(N303), .IN3(N304), .IN4(N305), .Q(n59) );
  NAND3X0 U577 ( .IN1(n1039), .IN2(n707), .IN3(N251), .QN(n67) );
  NAND3X0 U578 ( .IN1(n1036), .IN2(n1171), .IN3(tempA[31]), .QN(n66) );
  NAND3X0 U581 ( .IN1(n1039), .IN2(n1170), .IN3(tempA[31]), .QN(n73) );
  NAND3X0 U583 ( .IN1(n1036), .IN2(n707), .IN3(N285), .QN(n72) );
  AO222X1 U586 ( .IN1(tempB[31]), .IN2(n76), .IN3(n77), .IN4(n1033), .IN5(
        tempA[31]), .IN6(n1029), .Q(n75) );
  AO21X1 U588 ( .IN1(tempA[31]), .IN2(n1032), .IN3(n1027), .Q(n76) );
  AO222X1 U590 ( .IN1(tempB[30]), .IN2(n82), .IN3(n83), .IN4(n1035), .IN5(
        tempA[30]), .IN6(n1031), .Q(n81) );
  AO21X1 U592 ( .IN1(tempA[30]), .IN2(n80), .IN3(n1027), .Q(n82) );
  AO222X1 U594 ( .IN1(tempB[29]), .IN2(n85), .IN3(n86), .IN4(n1035), .IN5(
        tempA[29]), .IN6(n1031), .Q(n84) );
  AO21X1 U596 ( .IN1(tempA[29]), .IN2(n80), .IN3(n1027), .Q(n85) );
  AO222X1 U598 ( .IN1(tempB[28]), .IN2(n88), .IN3(n89), .IN4(n1035), .IN5(
        tempA[28]), .IN6(n1031), .Q(n87) );
  AO21X1 U600 ( .IN1(tempA[28]), .IN2(n80), .IN3(n1027), .Q(n88) );
  AO222X1 U602 ( .IN1(tempB[27]), .IN2(n91), .IN3(n92), .IN4(n1034), .IN5(
        tempA[27]), .IN6(n1031), .Q(n90) );
  AO21X1 U604 ( .IN1(tempA[27]), .IN2(n1032), .IN3(n1027), .Q(n91) );
  AO222X1 U606 ( .IN1(tempB[26]), .IN2(n94), .IN3(n95), .IN4(n1034), .IN5(
        tempA[26]), .IN6(n1031), .Q(n93) );
  AO21X1 U608 ( .IN1(tempA[26]), .IN2(n1032), .IN3(n1027), .Q(n94) );
  AO222X1 U610 ( .IN1(tempB[25]), .IN2(n97), .IN3(n98), .IN4(n1034), .IN5(
        tempA[25]), .IN6(n1031), .Q(n96) );
  AO21X1 U612 ( .IN1(tempA[25]), .IN2(n1032), .IN3(n1028), .Q(n97) );
  AO222X1 U614 ( .IN1(tempB[24]), .IN2(n100), .IN3(n101), .IN4(n1034), .IN5(
        tempA[24]), .IN6(n1031), .Q(n99) );
  AO21X1 U616 ( .IN1(tempA[24]), .IN2(n80), .IN3(n1028), .Q(n100) );
  AO222X1 U618 ( .IN1(tempB[23]), .IN2(n103), .IN3(n104), .IN4(n1034), .IN5(
        tempA[23]), .IN6(n1031), .Q(n102) );
  AO21X1 U620 ( .IN1(tempA[23]), .IN2(n1032), .IN3(n1028), .Q(n103) );
  AO222X1 U622 ( .IN1(tempB[22]), .IN2(n106), .IN3(n107), .IN4(n1034), .IN5(
        tempA[22]), .IN6(n1031), .Q(n105) );
  AO21X1 U624 ( .IN1(tempA[22]), .IN2(n1032), .IN3(n1028), .Q(n106) );
  AO222X1 U626 ( .IN1(tempB[21]), .IN2(n109), .IN3(n110), .IN4(n1034), .IN5(
        tempA[21]), .IN6(n1031), .Q(n108) );
  AO21X1 U628 ( .IN1(tempA[21]), .IN2(n1032), .IN3(n1028), .Q(n109) );
  AO222X1 U630 ( .IN1(tempB[20]), .IN2(n112), .IN3(n113), .IN4(n1034), .IN5(
        tempA[20]), .IN6(n1030), .Q(n111) );
  AO21X1 U632 ( .IN1(tempA[20]), .IN2(n1032), .IN3(n1028), .Q(n112) );
  AO222X1 U634 ( .IN1(tempB[19]), .IN2(n115), .IN3(n116), .IN4(n1034), .IN5(
        tempA[19]), .IN6(n1030), .Q(n114) );
  AO21X1 U636 ( .IN1(tempA[19]), .IN2(n1032), .IN3(n1028), .Q(n115) );
  AO222X1 U638 ( .IN1(tempB[18]), .IN2(n118), .IN3(n119), .IN4(n1034), .IN5(
        tempA[18]), .IN6(n1030), .Q(n117) );
  AO21X1 U640 ( .IN1(tempA[18]), .IN2(n1032), .IN3(n1028), .Q(n118) );
  AO222X1 U642 ( .IN1(tempB[17]), .IN2(n121), .IN3(n122), .IN4(n1034), .IN5(
        tempA[17]), .IN6(n1030), .Q(n120) );
  AO21X1 U644 ( .IN1(tempA[17]), .IN2(n1032), .IN3(n1028), .Q(n121) );
  AO222X1 U646 ( .IN1(tempB[16]), .IN2(n124), .IN3(n125), .IN4(n1034), .IN5(
        tempA[16]), .IN6(n1030), .Q(n123) );
  AO21X1 U648 ( .IN1(tempA[16]), .IN2(n1032), .IN3(n1029), .Q(n124) );
  AO222X1 U650 ( .IN1(tempB[15]), .IN2(n127), .IN3(n128), .IN4(n1034), .IN5(
        tempA[15]), .IN6(n1030), .Q(n126) );
  AO21X1 U652 ( .IN1(tempA[15]), .IN2(n1032), .IN3(n1029), .Q(n127) );
  AO222X1 U654 ( .IN1(tempB[14]), .IN2(n130), .IN3(n131), .IN4(n1034), .IN5(
        tempA[14]), .IN6(n1030), .Q(n129) );
  AO21X1 U656 ( .IN1(tempA[14]), .IN2(n1032), .IN3(n1029), .Q(n130) );
  AO222X1 U658 ( .IN1(tempB[13]), .IN2(n133), .IN3(n134), .IN4(n1033), .IN5(
        tempA[13]), .IN6(n1030), .Q(n132) );
  AO21X1 U660 ( .IN1(tempA[13]), .IN2(n80), .IN3(n1029), .Q(n133) );
  AO222X1 U662 ( .IN1(tempB[12]), .IN2(n136), .IN3(n137), .IN4(n1033), .IN5(
        tempA[12]), .IN6(n1030), .Q(n135) );
  AO21X1 U664 ( .IN1(tempA[12]), .IN2(n80), .IN3(n1029), .Q(n136) );
  AO222X1 U666 ( .IN1(tempB[11]), .IN2(n139), .IN3(n140), .IN4(n1033), .IN5(
        tempA[11]), .IN6(n1030), .Q(n138) );
  AO21X1 U668 ( .IN1(tempA[11]), .IN2(n1032), .IN3(n1028), .Q(n139) );
  AO222X1 U670 ( .IN1(tempB[10]), .IN2(n142), .IN3(n143), .IN4(n1033), .IN5(
        tempA[10]), .IN6(n1030), .Q(n141) );
  AO21X1 U672 ( .IN1(tempA[10]), .IN2(n1032), .IN3(n1029), .Q(n142) );
  AO222X1 U674 ( .IN1(tempB[9]), .IN2(n145), .IN3(n146), .IN4(n1033), .IN5(
        n1027), .IN6(tempA[9]), .Q(n144) );
  AO21X1 U676 ( .IN1(tempA[9]), .IN2(n1032), .IN3(n1027), .Q(n145) );
  AO222X1 U678 ( .IN1(tempB[8]), .IN2(n148), .IN3(n149), .IN4(n1033), .IN5(
        tempA[8]), .IN6(n1029), .Q(n147) );
  AO21X1 U680 ( .IN1(tempA[8]), .IN2(n1032), .IN3(n1028), .Q(n148) );
  AO222X1 U682 ( .IN1(tempB[7]), .IN2(n151), .IN3(n152), .IN4(n1034), .IN5(
        tempA[7]), .IN6(n1030), .Q(n150) );
  AO21X1 U684 ( .IN1(tempA[7]), .IN2(n1032), .IN3(n1028), .Q(n151) );
  AO222X1 U686 ( .IN1(tempB[6]), .IN2(n154), .IN3(n155), .IN4(n1033), .IN5(
        tempA[6]), .IN6(n1029), .Q(n153) );
  AO21X1 U688 ( .IN1(tempA[6]), .IN2(n1032), .IN3(n1027), .Q(n154) );
  AO222X1 U690 ( .IN1(tempB[5]), .IN2(n157), .IN3(n158), .IN4(n1033), .IN5(
        tempA[5]), .IN6(n1029), .Q(n156) );
  AO21X1 U692 ( .IN1(tempA[5]), .IN2(n1032), .IN3(n1028), .Q(n157) );
  AO222X1 U694 ( .IN1(tempB[4]), .IN2(n160), .IN3(n161), .IN4(n1033), .IN5(
        tempA[4]), .IN6(n1029), .Q(n159) );
  AO21X1 U696 ( .IN1(tempA[4]), .IN2(n1032), .IN3(n1027), .Q(n160) );
  AO222X1 U698 ( .IN1(tempB[3]), .IN2(n163), .IN3(n164), .IN4(n1033), .IN5(
        tempA[3]), .IN6(n1029), .Q(n162) );
  AO21X1 U700 ( .IN1(tempA[3]), .IN2(n1032), .IN3(n1027), .Q(n163) );
  AO222X1 U702 ( .IN1(tempB[2]), .IN2(n166), .IN3(n167), .IN4(n1033), .IN5(
        tempA[2]), .IN6(n1029), .Q(n165) );
  AO21X1 U704 ( .IN1(tempA[2]), .IN2(n1032), .IN3(n1027), .Q(n166) );
  AO222X1 U706 ( .IN1(tempB[1]), .IN2(n169), .IN3(n170), .IN4(n1033), .IN5(
        tempA[1]), .IN6(n1030), .Q(n168) );
  AO21X1 U708 ( .IN1(tempA[1]), .IN2(n1032), .IN3(n1027), .Q(n169) );
  AOI222X1 U710 ( .IN1(N254), .IN2(n1038), .IN3(tempA[0]), .IN4(n1031), .IN5(
        N220), .IN6(n1039), .QN(n174) );
  AO21X1 U712 ( .IN1(n175), .IN2(n176), .IN3(n705), .Q(n173) );
  NOR3X0 U715 ( .IN1(opcode[1]), .IN2(opcode[3]), .IN3(n702), .QN(n80) );
  NAND4X0 U716 ( .IN1(N288), .IN2(n179), .IN3(n183), .IN4(n702), .QN(n172) );
  NAND3X0 U717 ( .IN1(n710), .IN2(n705), .IN3(n1033), .QN(n171) );
  AO221X1 U720 ( .IN1(N252), .IN2(n1040), .IN3(N286), .IN4(n1037), .IN5(n1033), 
        .Q(N289) );
  AND4X1 U721 ( .IN1(opcode[3]), .IN2(n706), .IN3(n702), .IN4(n711), .Q(n78)
         );
  AND3X1 U722 ( .IN1(n706), .IN2(n702), .IN3(n179), .Q(n70) );
  AND3X1 U724 ( .IN1(n700), .IN2(n706), .IN3(n179), .Q(n68) );
  pipealu_DW_cmp_0 lt_73 ( .A(tempA), .B(tempB), .TC(1'b0), .GE_LT(1'b1), 
        .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N288) );
  pipealu_DW01_sub_0 sub_67 ( .A({1'b0, tempA}), .B({1'b0, tempB}), .CI(1'b0), 
        .DIFF({N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, 
        N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, 
        N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254}) );
  pipealu_DW01_add_0 add_61 ( .A({1'b0, tempA}), .B({1'b0, tempB}), .CI(1'b0), 
        .SUM({N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, 
        N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, 
        N229, N228, N227, N226, N225, N224, N223, N222, N221, N220}) );
  INVX0 U728 ( .INP(n1045), .ZN(n1043) );
  INVX0 U729 ( .INP(n1045), .ZN(n1042) );
  INVX0 U730 ( .INP(n52), .ZN(n1045) );
  INVX0 U731 ( .INP(n1141), .ZN(n1139) );
  INVX0 U732 ( .INP(n1109), .ZN(n1107) );
  INVX0 U733 ( .INP(n1085), .ZN(n1083) );
  INVX0 U734 ( .INP(n1117), .ZN(n1115) );
  INVX0 U735 ( .INP(n1149), .ZN(n1147) );
  INVX0 U736 ( .INP(n1157), .ZN(n1155) );
  INVX0 U737 ( .INP(n1053), .ZN(n1051) );
  INVX0 U738 ( .INP(n1061), .ZN(n1059) );
  INVX0 U739 ( .INP(n1093), .ZN(n1091) );
  INVX0 U740 ( .INP(n1101), .ZN(n1099) );
  INVX0 U741 ( .INP(n1133), .ZN(n1131) );
  INVX0 U742 ( .INP(n1165), .ZN(n1163) );
  INVX0 U743 ( .INP(n1077), .ZN(n1075) );
  INVX0 U744 ( .INP(n1125), .ZN(n1123) );
  INVX0 U745 ( .INP(n1069), .ZN(n1067) );
  INVX0 U746 ( .INP(n52), .ZN(n1049) );
  INVX0 U747 ( .INP(n52), .ZN(n1046) );
  INVX0 U748 ( .INP(n52), .ZN(n1047) );
  INVX0 U749 ( .INP(n52), .ZN(n1048) );
  INVX0 U750 ( .INP(n1141), .ZN(n1138) );
  INVX0 U751 ( .INP(n1109), .ZN(n1106) );
  INVX0 U752 ( .INP(n1085), .ZN(n1082) );
  INVX0 U753 ( .INP(n1117), .ZN(n1114) );
  INVX0 U754 ( .INP(n1149), .ZN(n1146) );
  INVX0 U755 ( .INP(n1157), .ZN(n1154) );
  INVX0 U756 ( .INP(n1053), .ZN(n1050) );
  INVX0 U757 ( .INP(n1061), .ZN(n1058) );
  INVX0 U758 ( .INP(n1093), .ZN(n1090) );
  INVX0 U759 ( .INP(n1101), .ZN(n1098) );
  INVX0 U760 ( .INP(n1133), .ZN(n1130) );
  INVX0 U761 ( .INP(n1165), .ZN(n1162) );
  INVX0 U762 ( .INP(n1077), .ZN(n1074) );
  INVX0 U763 ( .INP(n1125), .ZN(n1122) );
  INVX0 U764 ( .INP(n1069), .ZN(n1066) );
  NBUFFX2 U765 ( .INP(n70), .Z(n1038) );
  INVX0 U766 ( .INP(n46), .ZN(n1061) );
  INVX0 U767 ( .INP(n44), .ZN(n1069) );
  INVX0 U768 ( .INP(n41), .ZN(n1077) );
  INVX0 U769 ( .INP(n39), .ZN(n1085) );
  INVX0 U770 ( .INP(n36), .ZN(n1093) );
  INVX0 U771 ( .INP(n10), .ZN(n1165) );
  INVX0 U772 ( .INP(n26), .ZN(n1125) );
  INVX0 U773 ( .INP(n24), .ZN(n1133) );
  INVX0 U774 ( .INP(n17), .ZN(n1149) );
  INVX0 U775 ( .INP(n21), .ZN(n1141) );
  INVX0 U776 ( .INP(n48), .ZN(n1053) );
  INVX0 U777 ( .INP(n14), .ZN(n1157) );
  INVX0 U778 ( .INP(n34), .ZN(n1101) );
  INVX0 U779 ( .INP(n32), .ZN(n1109) );
  INVX0 U780 ( .INP(n29), .ZN(n1117) );
  NAND2X1 U781 ( .IN1(n30), .IN2(n15), .QN(n52) );
  INVX0 U782 ( .INP(n46), .ZN(n1065) );
  INVX0 U783 ( .INP(n46), .ZN(n1062) );
  INVX0 U784 ( .INP(n46), .ZN(n1063) );
  INVX0 U785 ( .INP(n46), .ZN(n1064) );
  INVX0 U786 ( .INP(n44), .ZN(n1073) );
  INVX0 U787 ( .INP(n44), .ZN(n1070) );
  INVX0 U788 ( .INP(n44), .ZN(n1071) );
  INVX0 U789 ( .INP(n44), .ZN(n1072) );
  INVX0 U790 ( .INP(n41), .ZN(n1081) );
  INVX0 U791 ( .INP(n41), .ZN(n1078) );
  INVX0 U792 ( .INP(n41), .ZN(n1079) );
  INVX0 U793 ( .INP(n41), .ZN(n1080) );
  INVX0 U794 ( .INP(n39), .ZN(n1089) );
  INVX0 U795 ( .INP(n39), .ZN(n1086) );
  INVX0 U796 ( .INP(n39), .ZN(n1087) );
  INVX0 U797 ( .INP(n39), .ZN(n1088) );
  INVX0 U798 ( .INP(n36), .ZN(n1097) );
  INVX0 U799 ( .INP(n36), .ZN(n1094) );
  INVX0 U800 ( .INP(n36), .ZN(n1095) );
  INVX0 U801 ( .INP(n36), .ZN(n1096) );
  INVX0 U802 ( .INP(n10), .ZN(n1169) );
  INVX0 U803 ( .INP(n10), .ZN(n1166) );
  INVX0 U804 ( .INP(n10), .ZN(n1167) );
  INVX0 U805 ( .INP(n10), .ZN(n1168) );
  INVX0 U806 ( .INP(n26), .ZN(n1129) );
  INVX0 U807 ( .INP(n26), .ZN(n1126) );
  INVX0 U808 ( .INP(n26), .ZN(n1127) );
  INVX0 U809 ( .INP(n26), .ZN(n1128) );
  INVX0 U810 ( .INP(n24), .ZN(n1137) );
  INVX0 U811 ( .INP(n24), .ZN(n1134) );
  INVX0 U812 ( .INP(n24), .ZN(n1135) );
  INVX0 U813 ( .INP(n24), .ZN(n1136) );
  INVX0 U814 ( .INP(n17), .ZN(n1153) );
  INVX0 U815 ( .INP(n17), .ZN(n1150) );
  INVX0 U816 ( .INP(n17), .ZN(n1151) );
  INVX0 U817 ( .INP(n17), .ZN(n1152) );
  INVX0 U818 ( .INP(n21), .ZN(n1145) );
  INVX0 U819 ( .INP(n21), .ZN(n1142) );
  INVX0 U820 ( .INP(n21), .ZN(n1143) );
  INVX0 U821 ( .INP(n21), .ZN(n1144) );
  INVX0 U822 ( .INP(n48), .ZN(n1057) );
  INVX0 U823 ( .INP(n48), .ZN(n1054) );
  INVX0 U824 ( .INP(n48), .ZN(n1055) );
  INVX0 U825 ( .INP(n48), .ZN(n1056) );
  INVX0 U826 ( .INP(n14), .ZN(n1161) );
  INVX0 U827 ( .INP(n14), .ZN(n1158) );
  INVX0 U828 ( .INP(n14), .ZN(n1159) );
  INVX0 U829 ( .INP(n14), .ZN(n1160) );
  INVX0 U830 ( .INP(n34), .ZN(n1105) );
  INVX0 U831 ( .INP(n34), .ZN(n1102) );
  INVX0 U832 ( .INP(n34), .ZN(n1103) );
  INVX0 U833 ( .INP(n34), .ZN(n1104) );
  INVX0 U834 ( .INP(n32), .ZN(n1113) );
  INVX0 U835 ( .INP(n32), .ZN(n1110) );
  INVX0 U836 ( .INP(n32), .ZN(n1111) );
  INVX0 U837 ( .INP(n32), .ZN(n1112) );
  INVX0 U838 ( .INP(n29), .ZN(n1121) );
  INVX0 U839 ( .INP(n29), .ZN(n1118) );
  INVX0 U840 ( .INP(n29), .ZN(n1119) );
  INVX0 U841 ( .INP(n29), .ZN(n1120) );
  INVX0 U842 ( .INP(n175), .ZN(n1172) );
  NOR2X0 U843 ( .IN1(n703), .IN2(n709), .QN(n15) );
  NOR2X0 U844 ( .IN1(n704), .IN2(n708), .QN(n30) );
  NAND2X1 U845 ( .IN1(n22), .IN2(n18), .QN(n21) );
  NAND2X1 U846 ( .IN1(n30), .IN2(n22), .QN(n32) );
  NAND2X1 U847 ( .IN1(n37), .IN2(n22), .QN(n39) );
  NAND2X1 U848 ( .IN1(n30), .IN2(n19), .QN(n29) );
  NAND2X1 U849 ( .IN1(n18), .IN2(n19), .QN(n17) );
  NAND2X1 U850 ( .IN1(n37), .IN2(n19), .QN(n36) );
  NAND2X1 U851 ( .IN1(n15), .IN2(n11), .QN(n14) );
  NAND2X1 U852 ( .IN1(n22), .IN2(n11), .QN(n48) );
  NAND2X1 U853 ( .IN1(n19), .IN2(n11), .QN(n46) );
  NAND2X1 U854 ( .IN1(n30), .IN2(n12), .QN(n34) );
  NAND2X1 U855 ( .IN1(n18), .IN2(n12), .QN(n24) );
  NAND2X1 U856 ( .IN1(n11), .IN2(n12), .QN(n10) );
  NAND2X1 U857 ( .IN1(n37), .IN2(n12), .QN(n41) );
  NAND2X1 U858 ( .IN1(n18), .IN2(n15), .QN(n26) );
  NAND2X1 U859 ( .IN1(n37), .IN2(n15), .QN(n44) );
  NBUFFX2 U860 ( .INP(n78), .Z(n1035) );
  NBUFFX2 U861 ( .INP(n68), .Z(n1041) );
  INVX0 U862 ( .INP(N251), .ZN(n1170) );
  AO221X1 U863 ( .IN1(N250), .IN2(n1041), .IN3(N284), .IN4(n1038), .IN5(n81), 
        .Q(N320) );
  NOR2X0 U864 ( .IN1(tempB[30]), .IN2(tempA[30]), .QN(n83) );
  AO221X1 U865 ( .IN1(N248), .IN2(n1040), .IN3(N282), .IN4(n1038), .IN5(n87), 
        .Q(N318) );
  NOR2X0 U866 ( .IN1(tempB[28]), .IN2(tempA[28]), .QN(n89) );
  AO221X1 U867 ( .IN1(N249), .IN2(n1041), .IN3(N283), .IN4(n1038), .IN5(n84), 
        .Q(N319) );
  NOR2X0 U868 ( .IN1(tempB[29]), .IN2(tempA[29]), .QN(n86) );
  AO221X1 U869 ( .IN1(N246), .IN2(n1040), .IN3(N280), .IN4(n1038), .IN5(n93), 
        .Q(N316) );
  NOR2X0 U870 ( .IN1(tempB[26]), .IN2(tempA[26]), .QN(n95) );
  AO221X1 U871 ( .IN1(N245), .IN2(n1040), .IN3(N279), .IN4(n1037), .IN5(n96), 
        .Q(N315) );
  NOR2X0 U872 ( .IN1(tempB[25]), .IN2(tempA[25]), .QN(n98) );
  AO221X1 U873 ( .IN1(N247), .IN2(n1040), .IN3(N281), .IN4(n1038), .IN5(n90), 
        .Q(N317) );
  NOR2X0 U874 ( .IN1(tempB[27]), .IN2(tempA[27]), .QN(n92) );
  AO221X1 U875 ( .IN1(N251), .IN2(n1039), .IN3(N285), .IN4(n1036), .IN5(n75), 
        .Q(N321) );
  NOR2X0 U876 ( .IN1(tempB[31]), .IN2(tempA[31]), .QN(n77) );
  OAI22X1 U877 ( .IN1(n712), .IN2(n713), .IN3(n714), .IN4(tempB[31]), .QN(N322) );
  AND2X1 U878 ( .IN1(n72), .IN2(n73), .Q(n713) );
  AND2X1 U879 ( .IN1(n66), .IN2(n67), .Q(n714) );
  INVX0 U880 ( .INP(N285), .ZN(n1171) );
  AO221X1 U881 ( .IN1(N236), .IN2(n1040), .IN3(N270), .IN4(n1037), .IN5(n123), 
        .Q(N306) );
  NOR2X0 U882 ( .IN1(tempB[16]), .IN2(tempA[16]), .QN(n125) );
  AO221X1 U883 ( .IN1(N240), .IN2(n1040), .IN3(N274), .IN4(n1037), .IN5(n111), 
        .Q(N310) );
  NOR2X0 U884 ( .IN1(tempB[20]), .IN2(tempA[20]), .QN(n113) );
  AO221X1 U885 ( .IN1(N244), .IN2(n1040), .IN3(N278), .IN4(n1037), .IN5(n99), 
        .Q(N314) );
  NOR2X0 U886 ( .IN1(tempB[24]), .IN2(tempA[24]), .QN(n101) );
  AO221X1 U887 ( .IN1(N234), .IN2(n1040), .IN3(N268), .IN4(n1037), .IN5(n129), 
        .Q(N304) );
  NOR2X0 U888 ( .IN1(tempB[14]), .IN2(tempA[14]), .QN(n131) );
  AO221X1 U889 ( .IN1(N238), .IN2(n1040), .IN3(N272), .IN4(n1037), .IN5(n117), 
        .Q(N308) );
  NOR2X0 U890 ( .IN1(tempB[18]), .IN2(tempA[18]), .QN(n119) );
  AO221X1 U891 ( .IN1(N242), .IN2(n1040), .IN3(N276), .IN4(n1037), .IN5(n105), 
        .Q(N312) );
  NOR2X0 U892 ( .IN1(tempB[22]), .IN2(tempA[22]), .QN(n107) );
  AO221X1 U893 ( .IN1(N237), .IN2(n1040), .IN3(N271), .IN4(n1037), .IN5(n120), 
        .Q(N307) );
  NOR2X0 U894 ( .IN1(tempB[17]), .IN2(tempA[17]), .QN(n122) );
  AO221X1 U895 ( .IN1(N241), .IN2(n1040), .IN3(N275), .IN4(n1037), .IN5(n108), 
        .Q(N311) );
  NOR2X0 U896 ( .IN1(tempB[21]), .IN2(tempA[21]), .QN(n110) );
  AO221X1 U897 ( .IN1(N235), .IN2(n1040), .IN3(N269), .IN4(n1037), .IN5(n126), 
        .Q(N305) );
  NOR2X0 U898 ( .IN1(tempB[15]), .IN2(tempA[15]), .QN(n128) );
  AO221X1 U899 ( .IN1(N239), .IN2(n1040), .IN3(N273), .IN4(n1037), .IN5(n114), 
        .Q(N309) );
  NOR2X0 U900 ( .IN1(tempB[19]), .IN2(tempA[19]), .QN(n116) );
  AO221X1 U901 ( .IN1(N243), .IN2(n1040), .IN3(N277), .IN4(n1037), .IN5(n102), 
        .Q(N313) );
  NOR2X0 U902 ( .IN1(tempB[23]), .IN2(tempA[23]), .QN(n104) );
  NAND4X0 U903 ( .IN1(n171), .IN2(n172), .IN3(n173), .IN4(n174), .QN(N290) );
  AO221X1 U904 ( .IN1(N228), .IN2(n1039), .IN3(N262), .IN4(n1036), .IN5(n147), 
        .Q(N298) );
  NOR2X0 U905 ( .IN1(tempB[8]), .IN2(tempA[8]), .QN(n149) );
  AO221X1 U906 ( .IN1(N232), .IN2(n1039), .IN3(N266), .IN4(n1037), .IN5(n135), 
        .Q(N302) );
  NOR2X0 U907 ( .IN1(tempB[12]), .IN2(tempA[12]), .QN(n137) );
  AO221X1 U908 ( .IN1(N230), .IN2(n1039), .IN3(N264), .IN4(n1036), .IN5(n141), 
        .Q(N300) );
  NOR2X0 U909 ( .IN1(tempB[10]), .IN2(tempA[10]), .QN(n143) );
  AO221X1 U910 ( .IN1(N229), .IN2(n1039), .IN3(N263), .IN4(n1036), .IN5(n144), 
        .Q(N299) );
  NOR2X0 U911 ( .IN1(tempB[9]), .IN2(tempA[9]), .QN(n146) );
  AO221X1 U912 ( .IN1(N233), .IN2(n1040), .IN3(N267), .IN4(n1037), .IN5(n132), 
        .Q(N303) );
  NOR2X0 U913 ( .IN1(tempB[13]), .IN2(tempA[13]), .QN(n134) );
  AO221X1 U914 ( .IN1(N227), .IN2(n1039), .IN3(N261), .IN4(n1036), .IN5(n150), 
        .Q(N297) );
  NOR2X0 U915 ( .IN1(tempB[7]), .IN2(tempA[7]), .QN(n152) );
  AO221X1 U916 ( .IN1(N231), .IN2(n1039), .IN3(N265), .IN4(n1036), .IN5(n138), 
        .Q(N301) );
  NOR2X0 U917 ( .IN1(tempB[11]), .IN2(tempA[11]), .QN(n140) );
  NAND2X1 U918 ( .IN1(n183), .IN2(n1032), .QN(n175) );
  NAND2X1 U919 ( .IN1(tempA[0]), .IN2(n80), .QN(n176) );
  AO221X1 U920 ( .IN1(N221), .IN2(n1039), .IN3(N255), .IN4(n1036), .IN5(n168), 
        .Q(N291) );
  NOR2X0 U921 ( .IN1(tempB[1]), .IN2(tempA[1]), .QN(n170) );
  AO221X1 U922 ( .IN1(N223), .IN2(n1039), .IN3(N257), .IN4(n1036), .IN5(n162), 
        .Q(N293) );
  NOR2X0 U923 ( .IN1(tempB[3]), .IN2(tempA[3]), .QN(n164) );
  AO221X1 U924 ( .IN1(N224), .IN2(n1039), .IN3(N258), .IN4(n1036), .IN5(n159), 
        .Q(N294) );
  NOR2X0 U925 ( .IN1(tempB[4]), .IN2(tempA[4]), .QN(n161) );
  AO221X1 U926 ( .IN1(N225), .IN2(n1039), .IN3(N259), .IN4(n1036), .IN5(n156), 
        .Q(N295) );
  NOR2X0 U927 ( .IN1(tempB[5]), .IN2(tempA[5]), .QN(n158) );
  AO221X1 U928 ( .IN1(N222), .IN2(n1039), .IN3(N256), .IN4(n1036), .IN5(n165), 
        .Q(N292) );
  NOR2X0 U929 ( .IN1(tempB[2]), .IN2(tempA[2]), .QN(n167) );
  AO221X1 U930 ( .IN1(N226), .IN2(n1039), .IN3(N260), .IN4(n1036), .IN5(n153), 
        .Q(N296) );
  NOR2X0 U931 ( .IN1(tempB[6]), .IN2(tempA[6]), .QN(n155) );
  NOR2X0 U932 ( .IN1(n711), .IN2(opcode[3]), .QN(n179) );
  NOR2X0 U933 ( .IN1(n187), .IN2(n186), .QN(n19) );
  NOR2X0 U934 ( .IN1(n185), .IN2(n184), .QN(n37) );
  NOR2X0 U935 ( .IN1(n709), .IN2(n186), .QN(n12) );
  NOR2X0 U936 ( .IN1(n708), .IN2(n185), .QN(n11) );
  NOR2X0 U937 ( .IN1(n704), .IN2(n184), .QN(n18) );
  NOR2X0 U938 ( .IN1(n703), .IN2(n187), .QN(n22) );
  NBUFFX2 U939 ( .INP(N18), .Z(n854) );
  NBUFFX2 U940 ( .INP(N22), .Z(n1010) );
  NBUFFX2 U941 ( .INP(N17), .Z(n843) );
  NBUFFX2 U942 ( .INP(N21), .Z(n999) );
  NBUFFX2 U943 ( .INP(N19), .Z(n865) );
  NBUFFX2 U944 ( .INP(N23), .Z(n1021) );
  NBUFFX4 U945 ( .INP(N17), .Z(n844) );
  NBUFFX4 U946 ( .INP(N17), .Z(n845) );
  NBUFFX4 U947 ( .INP(N17), .Z(n846) );
  NBUFFX4 U948 ( .INP(N17), .Z(n847) );
  NBUFFX4 U949 ( .INP(N17), .Z(n848) );
  NBUFFX4 U950 ( .INP(N17), .Z(n849) );
  NBUFFX4 U951 ( .INP(N17), .Z(n850) );
  NBUFFX4 U952 ( .INP(N17), .Z(n851) );
  NBUFFX4 U953 ( .INP(N17), .Z(n852) );
  NBUFFX4 U954 ( .INP(N17), .Z(n853) );
  NBUFFX4 U955 ( .INP(N21), .Z(n1000) );
  NBUFFX4 U956 ( .INP(N21), .Z(n1001) );
  NBUFFX4 U957 ( .INP(N21), .Z(n1002) );
  NBUFFX4 U958 ( .INP(N21), .Z(n1003) );
  NBUFFX4 U959 ( .INP(N21), .Z(n1004) );
  NBUFFX4 U960 ( .INP(N21), .Z(n1005) );
  NBUFFX4 U961 ( .INP(N21), .Z(n1006) );
  NBUFFX4 U962 ( .INP(N21), .Z(n1007) );
  NBUFFX4 U963 ( .INP(N21), .Z(n1008) );
  NBUFFX4 U964 ( .INP(N21), .Z(n1009) );
  NBUFFX4 U965 ( .INP(N19), .Z(n866) );
  NBUFFX4 U966 ( .INP(N19), .Z(n867) );
  NBUFFX4 U967 ( .INP(N23), .Z(n1022) );
  NBUFFX4 U968 ( .INP(N23), .Z(n1023) );
  NBUFFX2 U969 ( .INP(N20), .Z(n868) );
  NBUFFX2 U970 ( .INP(N24), .Z(n1024) );
  MUX41X1 U971 ( .IN1(\regfile[12][0] ), .IN3(\regfile[14][0] ), .IN2(
        \regfile[13][0] ), .IN4(\regfile[15][0] ), .S0(n854), .S1(n843), .Q(
        n715) );
  MUX41X1 U972 ( .IN1(\regfile[8][0] ), .IN3(\regfile[10][0] ), .IN2(
        \regfile[9][0] ), .IN4(\regfile[11][0] ), .S0(n854), .S1(n843), .Q(
        n716) );
  MUX41X1 U973 ( .IN1(\regfile[4][0] ), .IN3(\regfile[6][0] ), .IN2(
        \regfile[5][0] ), .IN4(\regfile[7][0] ), .S0(n854), .S1(n843), .Q(n717) );
  MUX41X1 U974 ( .IN1(\regfile[0][0] ), .IN3(\regfile[2][0] ), .IN2(
        \regfile[1][0] ), .IN4(\regfile[3][0] ), .S0(n854), .S1(n843), .Q(n718) );
  MUX41X1 U975 ( .IN1(n718), .IN3(n716), .IN2(n717), .IN4(n715), .S0(n868), 
        .S1(n865), .Q(N56) );
  MUX41X1 U976 ( .IN1(\regfile[12][1] ), .IN3(\regfile[14][1] ), .IN2(
        \regfile[13][1] ), .IN4(\regfile[15][1] ), .S0(n854), .S1(n843), .Q(
        n719) );
  MUX41X1 U977 ( .IN1(\regfile[8][1] ), .IN3(\regfile[10][1] ), .IN2(
        \regfile[9][1] ), .IN4(\regfile[11][1] ), .S0(n854), .S1(n843), .Q(
        n720) );
  MUX41X1 U978 ( .IN1(\regfile[4][1] ), .IN3(\regfile[6][1] ), .IN2(
        \regfile[5][1] ), .IN4(\regfile[7][1] ), .S0(n854), .S1(n843), .Q(n721) );
  MUX41X1 U979 ( .IN1(\regfile[0][1] ), .IN3(\regfile[2][1] ), .IN2(
        \regfile[1][1] ), .IN4(\regfile[3][1] ), .S0(n854), .S1(n843), .Q(n722) );
  MUX41X1 U980 ( .IN1(n722), .IN3(n720), .IN2(n721), .IN4(n719), .S0(n868), 
        .S1(n865), .Q(N55) );
  MUX41X1 U981 ( .IN1(\regfile[12][2] ), .IN3(\regfile[14][2] ), .IN2(
        \regfile[13][2] ), .IN4(\regfile[15][2] ), .S0(n855), .S1(n844), .Q(
        n723) );
  MUX41X1 U982 ( .IN1(\regfile[8][2] ), .IN3(\regfile[10][2] ), .IN2(
        \regfile[9][2] ), .IN4(\regfile[11][2] ), .S0(n855), .S1(n844), .Q(
        n724) );
  MUX41X1 U983 ( .IN1(\regfile[4][2] ), .IN3(\regfile[6][2] ), .IN2(
        \regfile[5][2] ), .IN4(\regfile[7][2] ), .S0(n855), .S1(n844), .Q(n725) );
  MUX41X1 U984 ( .IN1(\regfile[0][2] ), .IN3(\regfile[2][2] ), .IN2(
        \regfile[1][2] ), .IN4(\regfile[3][2] ), .S0(n855), .S1(n844), .Q(n726) );
  MUX41X1 U985 ( .IN1(n726), .IN3(n724), .IN2(n725), .IN4(n723), .S0(n868), 
        .S1(n865), .Q(N54) );
  MUX41X1 U986 ( .IN1(\regfile[12][3] ), .IN3(\regfile[14][3] ), .IN2(
        \regfile[13][3] ), .IN4(\regfile[15][3] ), .S0(n855), .S1(n844), .Q(
        n727) );
  MUX41X1 U987 ( .IN1(\regfile[8][3] ), .IN3(\regfile[10][3] ), .IN2(
        \regfile[9][3] ), .IN4(\regfile[11][3] ), .S0(n855), .S1(n844), .Q(
        n728) );
  MUX41X1 U988 ( .IN1(\regfile[4][3] ), .IN3(\regfile[6][3] ), .IN2(
        \regfile[5][3] ), .IN4(\regfile[7][3] ), .S0(n855), .S1(n844), .Q(n729) );
  MUX41X1 U989 ( .IN1(\regfile[0][3] ), .IN3(\regfile[2][3] ), .IN2(
        \regfile[1][3] ), .IN4(\regfile[3][3] ), .S0(n855), .S1(n844), .Q(n730) );
  MUX41X1 U990 ( .IN1(n730), .IN3(n728), .IN2(n729), .IN4(n727), .S0(n868), 
        .S1(n865), .Q(N53) );
  MUX41X1 U991 ( .IN1(\regfile[12][4] ), .IN3(\regfile[14][4] ), .IN2(
        \regfile[13][4] ), .IN4(\regfile[15][4] ), .S0(n855), .S1(n844), .Q(
        n731) );
  MUX41X1 U992 ( .IN1(\regfile[8][4] ), .IN3(\regfile[10][4] ), .IN2(
        \regfile[9][4] ), .IN4(\regfile[11][4] ), .S0(n855), .S1(n844), .Q(
        n732) );
  MUX41X1 U993 ( .IN1(\regfile[4][4] ), .IN3(\regfile[6][4] ), .IN2(
        \regfile[5][4] ), .IN4(\regfile[7][4] ), .S0(n855), .S1(n844), .Q(n733) );
  MUX41X1 U994 ( .IN1(\regfile[0][4] ), .IN3(\regfile[2][4] ), .IN2(
        \regfile[1][4] ), .IN4(\regfile[3][4] ), .S0(n855), .S1(n844), .Q(n734) );
  MUX41X1 U995 ( .IN1(n734), .IN3(n732), .IN2(n733), .IN4(n731), .S0(n868), 
        .S1(n865), .Q(N52) );
  MUX41X1 U996 ( .IN1(\regfile[12][5] ), .IN3(\regfile[14][5] ), .IN2(
        \regfile[13][5] ), .IN4(\regfile[15][5] ), .S0(n856), .S1(n845), .Q(
        n735) );
  MUX41X1 U997 ( .IN1(\regfile[8][5] ), .IN3(\regfile[10][5] ), .IN2(
        \regfile[9][5] ), .IN4(\regfile[11][5] ), .S0(n856), .S1(n845), .Q(
        n736) );
  MUX41X1 U998 ( .IN1(\regfile[4][5] ), .IN3(\regfile[6][5] ), .IN2(
        \regfile[5][5] ), .IN4(\regfile[7][5] ), .S0(n856), .S1(n845), .Q(n737) );
  MUX41X1 U999 ( .IN1(\regfile[0][5] ), .IN3(\regfile[2][5] ), .IN2(
        \regfile[1][5] ), .IN4(\regfile[3][5] ), .S0(n856), .S1(n845), .Q(n738) );
  MUX41X1 U1000 ( .IN1(n738), .IN3(n736), .IN2(n737), .IN4(n735), .S0(n868), 
        .S1(n865), .Q(N51) );
  MUX41X1 U1001 ( .IN1(\regfile[12][6] ), .IN3(\regfile[14][6] ), .IN2(
        \regfile[13][6] ), .IN4(\regfile[15][6] ), .S0(n856), .S1(n845), .Q(
        n739) );
  MUX41X1 U1002 ( .IN1(\regfile[8][6] ), .IN3(\regfile[10][6] ), .IN2(
        \regfile[9][6] ), .IN4(\regfile[11][6] ), .S0(n856), .S1(n845), .Q(
        n740) );
  MUX41X1 U1003 ( .IN1(\regfile[4][6] ), .IN3(\regfile[6][6] ), .IN2(
        \regfile[5][6] ), .IN4(\regfile[7][6] ), .S0(n856), .S1(n845), .Q(n741) );
  MUX41X1 U1004 ( .IN1(\regfile[0][6] ), .IN3(\regfile[2][6] ), .IN2(
        \regfile[1][6] ), .IN4(\regfile[3][6] ), .S0(n856), .S1(n845), .Q(n742) );
  MUX41X1 U1005 ( .IN1(n742), .IN3(n740), .IN2(n741), .IN4(n739), .S0(n868), 
        .S1(n865), .Q(N50) );
  MUX41X1 U1006 ( .IN1(\regfile[12][7] ), .IN3(\regfile[14][7] ), .IN2(
        \regfile[13][7] ), .IN4(\regfile[15][7] ), .S0(n856), .S1(n845), .Q(
        n743) );
  MUX41X1 U1007 ( .IN1(\regfile[8][7] ), .IN3(\regfile[10][7] ), .IN2(
        \regfile[9][7] ), .IN4(\regfile[11][7] ), .S0(n856), .S1(n845), .Q(
        n744) );
  MUX41X1 U1008 ( .IN1(\regfile[4][7] ), .IN3(\regfile[6][7] ), .IN2(
        \regfile[5][7] ), .IN4(\regfile[7][7] ), .S0(n856), .S1(n845), .Q(n745) );
  MUX41X1 U1009 ( .IN1(\regfile[0][7] ), .IN3(\regfile[2][7] ), .IN2(
        \regfile[1][7] ), .IN4(\regfile[3][7] ), .S0(n856), .S1(n845), .Q(n746) );
  MUX41X1 U1010 ( .IN1(n746), .IN3(n744), .IN2(n745), .IN4(n743), .S0(n868), 
        .S1(n865), .Q(N49) );
  MUX41X1 U1011 ( .IN1(\regfile[12][8] ), .IN3(\regfile[14][8] ), .IN2(
        \regfile[13][8] ), .IN4(\regfile[15][8] ), .S0(n857), .S1(n846), .Q(
        n747) );
  MUX41X1 U1012 ( .IN1(\regfile[8][8] ), .IN3(\regfile[10][8] ), .IN2(
        \regfile[9][8] ), .IN4(\regfile[11][8] ), .S0(n857), .S1(n846), .Q(
        n748) );
  MUX41X1 U1013 ( .IN1(\regfile[4][8] ), .IN3(\regfile[6][8] ), .IN2(
        \regfile[5][8] ), .IN4(\regfile[7][8] ), .S0(n857), .S1(n846), .Q(n749) );
  MUX41X1 U1014 ( .IN1(\regfile[0][8] ), .IN3(\regfile[2][8] ), .IN2(
        \regfile[1][8] ), .IN4(\regfile[3][8] ), .S0(n857), .S1(n846), .Q(n750) );
  MUX41X1 U1015 ( .IN1(n750), .IN3(n748), .IN2(n749), .IN4(n747), .S0(n869), 
        .S1(n866), .Q(N48) );
  MUX41X1 U1016 ( .IN1(\regfile[12][9] ), .IN3(\regfile[14][9] ), .IN2(
        \regfile[13][9] ), .IN4(\regfile[15][9] ), .S0(n857), .S1(n846), .Q(
        n751) );
  MUX41X1 U1017 ( .IN1(\regfile[8][9] ), .IN3(\regfile[10][9] ), .IN2(
        \regfile[9][9] ), .IN4(\regfile[11][9] ), .S0(n857), .S1(n846), .Q(
        n752) );
  MUX41X1 U1018 ( .IN1(\regfile[4][9] ), .IN3(\regfile[6][9] ), .IN2(
        \regfile[5][9] ), .IN4(\regfile[7][9] ), .S0(n857), .S1(n846), .Q(n753) );
  MUX41X1 U1019 ( .IN1(\regfile[0][9] ), .IN3(\regfile[2][9] ), .IN2(
        \regfile[1][9] ), .IN4(\regfile[3][9] ), .S0(n857), .S1(n846), .Q(n754) );
  MUX41X1 U1020 ( .IN1(n754), .IN3(n752), .IN2(n753), .IN4(n751), .S0(n869), 
        .S1(n866), .Q(N47) );
  MUX41X1 U1021 ( .IN1(\regfile[12][10] ), .IN3(\regfile[14][10] ), .IN2(
        \regfile[13][10] ), .IN4(\regfile[15][10] ), .S0(n857), .S1(n846), .Q(
        n755) );
  MUX41X1 U1022 ( .IN1(\regfile[8][10] ), .IN3(\regfile[10][10] ), .IN2(
        \regfile[9][10] ), .IN4(\regfile[11][10] ), .S0(n857), .S1(n846), .Q(
        n756) );
  MUX41X1 U1023 ( .IN1(\regfile[4][10] ), .IN3(\regfile[6][10] ), .IN2(
        \regfile[5][10] ), .IN4(\regfile[7][10] ), .S0(n857), .S1(n846), .Q(
        n757) );
  MUX41X1 U1024 ( .IN1(\regfile[0][10] ), .IN3(\regfile[2][10] ), .IN2(
        \regfile[1][10] ), .IN4(\regfile[3][10] ), .S0(n857), .S1(n846), .Q(
        n758) );
  MUX41X1 U1025 ( .IN1(n758), .IN3(n756), .IN2(n757), .IN4(n755), .S0(n869), 
        .S1(n866), .Q(N46) );
  MUX41X1 U1026 ( .IN1(\regfile[12][11] ), .IN3(\regfile[14][11] ), .IN2(
        \regfile[13][11] ), .IN4(\regfile[15][11] ), .S0(n858), .S1(n847), .Q(
        n759) );
  MUX41X1 U1027 ( .IN1(\regfile[8][11] ), .IN3(\regfile[10][11] ), .IN2(
        \regfile[9][11] ), .IN4(\regfile[11][11] ), .S0(n858), .S1(n847), .Q(
        n760) );
  MUX41X1 U1028 ( .IN1(\regfile[4][11] ), .IN3(\regfile[6][11] ), .IN2(
        \regfile[5][11] ), .IN4(\regfile[7][11] ), .S0(n858), .S1(n847), .Q(
        n761) );
  MUX41X1 U1029 ( .IN1(\regfile[0][11] ), .IN3(\regfile[2][11] ), .IN2(
        \regfile[1][11] ), .IN4(\regfile[3][11] ), .S0(n858), .S1(n847), .Q(
        n762) );
  MUX41X1 U1030 ( .IN1(n762), .IN3(n760), .IN2(n761), .IN4(n759), .S0(n869), 
        .S1(n866), .Q(N45) );
  MUX41X1 U1031 ( .IN1(\regfile[12][12] ), .IN3(\regfile[14][12] ), .IN2(
        \regfile[13][12] ), .IN4(\regfile[15][12] ), .S0(n858), .S1(n847), .Q(
        n763) );
  MUX41X1 U1032 ( .IN1(\regfile[8][12] ), .IN3(\regfile[10][12] ), .IN2(
        \regfile[9][12] ), .IN4(\regfile[11][12] ), .S0(n858), .S1(n847), .Q(
        n764) );
  MUX41X1 U1033 ( .IN1(\regfile[4][12] ), .IN3(\regfile[6][12] ), .IN2(
        \regfile[5][12] ), .IN4(\regfile[7][12] ), .S0(n858), .S1(n847), .Q(
        n765) );
  MUX41X1 U1034 ( .IN1(\regfile[0][12] ), .IN3(\regfile[2][12] ), .IN2(
        \regfile[1][12] ), .IN4(\regfile[3][12] ), .S0(n858), .S1(n847), .Q(
        n766) );
  MUX41X1 U1035 ( .IN1(n766), .IN3(n764), .IN2(n765), .IN4(n763), .S0(n869), 
        .S1(n866), .Q(N44) );
  MUX41X1 U1036 ( .IN1(\regfile[12][13] ), .IN3(\regfile[14][13] ), .IN2(
        \regfile[13][13] ), .IN4(\regfile[15][13] ), .S0(n858), .S1(n847), .Q(
        n767) );
  MUX41X1 U1037 ( .IN1(\regfile[8][13] ), .IN3(\regfile[10][13] ), .IN2(
        \regfile[9][13] ), .IN4(\regfile[11][13] ), .S0(n858), .S1(n847), .Q(
        n768) );
  MUX41X1 U1038 ( .IN1(\regfile[4][13] ), .IN3(\regfile[6][13] ), .IN2(
        \regfile[5][13] ), .IN4(\regfile[7][13] ), .S0(n858), .S1(n847), .Q(
        n769) );
  MUX41X1 U1039 ( .IN1(\regfile[0][13] ), .IN3(\regfile[2][13] ), .IN2(
        \regfile[1][13] ), .IN4(\regfile[3][13] ), .S0(n858), .S1(n847), .Q(
        n770) );
  MUX41X1 U1040 ( .IN1(n770), .IN3(n768), .IN2(n769), .IN4(n767), .S0(n869), 
        .S1(n866), .Q(N43) );
  MUX41X1 U1041 ( .IN1(\regfile[12][14] ), .IN3(\regfile[14][14] ), .IN2(
        \regfile[13][14] ), .IN4(\regfile[15][14] ), .S0(n859), .S1(n848), .Q(
        n771) );
  MUX41X1 U1042 ( .IN1(\regfile[8][14] ), .IN3(\regfile[10][14] ), .IN2(
        \regfile[9][14] ), .IN4(\regfile[11][14] ), .S0(n859), .S1(n848), .Q(
        n772) );
  MUX41X1 U1043 ( .IN1(\regfile[4][14] ), .IN3(\regfile[6][14] ), .IN2(
        \regfile[5][14] ), .IN4(\regfile[7][14] ), .S0(n859), .S1(n848), .Q(
        n773) );
  MUX41X1 U1044 ( .IN1(\regfile[0][14] ), .IN3(\regfile[2][14] ), .IN2(
        \regfile[1][14] ), .IN4(\regfile[3][14] ), .S0(n859), .S1(n848), .Q(
        n774) );
  MUX41X1 U1045 ( .IN1(n774), .IN3(n772), .IN2(n773), .IN4(n771), .S0(n869), 
        .S1(n866), .Q(N42) );
  MUX41X1 U1046 ( .IN1(\regfile[12][15] ), .IN3(\regfile[14][15] ), .IN2(
        \regfile[13][15] ), .IN4(\regfile[15][15] ), .S0(n859), .S1(n848), .Q(
        n775) );
  MUX41X1 U1047 ( .IN1(\regfile[8][15] ), .IN3(\regfile[10][15] ), .IN2(
        \regfile[9][15] ), .IN4(\regfile[11][15] ), .S0(n859), .S1(n848), .Q(
        n776) );
  MUX41X1 U1048 ( .IN1(\regfile[4][15] ), .IN3(\regfile[6][15] ), .IN2(
        \regfile[5][15] ), .IN4(\regfile[7][15] ), .S0(n859), .S1(n848), .Q(
        n777) );
  MUX41X1 U1049 ( .IN1(\regfile[0][15] ), .IN3(\regfile[2][15] ), .IN2(
        \regfile[1][15] ), .IN4(\regfile[3][15] ), .S0(n859), .S1(n848), .Q(
        n778) );
  MUX41X1 U1050 ( .IN1(n778), .IN3(n776), .IN2(n777), .IN4(n775), .S0(n869), 
        .S1(n866), .Q(N41) );
  MUX41X1 U1051 ( .IN1(\regfile[12][16] ), .IN3(\regfile[14][16] ), .IN2(
        \regfile[13][16] ), .IN4(\regfile[15][16] ), .S0(n859), .S1(n848), .Q(
        n779) );
  MUX41X1 U1052 ( .IN1(\regfile[8][16] ), .IN3(\regfile[10][16] ), .IN2(
        \regfile[9][16] ), .IN4(\regfile[11][16] ), .S0(n859), .S1(n848), .Q(
        n780) );
  MUX41X1 U1053 ( .IN1(\regfile[4][16] ), .IN3(\regfile[6][16] ), .IN2(
        \regfile[5][16] ), .IN4(\regfile[7][16] ), .S0(n859), .S1(n848), .Q(
        n781) );
  MUX41X1 U1054 ( .IN1(\regfile[0][16] ), .IN3(\regfile[2][16] ), .IN2(
        \regfile[1][16] ), .IN4(\regfile[3][16] ), .S0(n859), .S1(n848), .Q(
        n782) );
  MUX41X1 U1055 ( .IN1(n782), .IN3(n780), .IN2(n781), .IN4(n779), .S0(n869), 
        .S1(n866), .Q(N40) );
  MUX41X1 U1056 ( .IN1(\regfile[12][17] ), .IN3(\regfile[14][17] ), .IN2(
        \regfile[13][17] ), .IN4(\regfile[15][17] ), .S0(n860), .S1(n849), .Q(
        n783) );
  MUX41X1 U1057 ( .IN1(\regfile[8][17] ), .IN3(\regfile[10][17] ), .IN2(
        \regfile[9][17] ), .IN4(\regfile[11][17] ), .S0(n860), .S1(n849), .Q(
        n784) );
  MUX41X1 U1058 ( .IN1(\regfile[4][17] ), .IN3(\regfile[6][17] ), .IN2(
        \regfile[5][17] ), .IN4(\regfile[7][17] ), .S0(n860), .S1(n849), .Q(
        n785) );
  MUX41X1 U1059 ( .IN1(\regfile[0][17] ), .IN3(\regfile[2][17] ), .IN2(
        \regfile[1][17] ), .IN4(\regfile[3][17] ), .S0(n860), .S1(n849), .Q(
        n786) );
  MUX41X1 U1060 ( .IN1(n786), .IN3(n784), .IN2(n785), .IN4(n783), .S0(n869), 
        .S1(n866), .Q(N39) );
  MUX41X1 U1061 ( .IN1(\regfile[12][18] ), .IN3(\regfile[14][18] ), .IN2(
        \regfile[13][18] ), .IN4(\regfile[15][18] ), .S0(n860), .S1(n849), .Q(
        n787) );
  MUX41X1 U1062 ( .IN1(\regfile[8][18] ), .IN3(\regfile[10][18] ), .IN2(
        \regfile[9][18] ), .IN4(\regfile[11][18] ), .S0(n860), .S1(n849), .Q(
        n788) );
  MUX41X1 U1063 ( .IN1(\regfile[4][18] ), .IN3(\regfile[6][18] ), .IN2(
        \regfile[5][18] ), .IN4(\regfile[7][18] ), .S0(n860), .S1(n849), .Q(
        n789) );
  MUX41X1 U1064 ( .IN1(\regfile[0][18] ), .IN3(\regfile[2][18] ), .IN2(
        \regfile[1][18] ), .IN4(\regfile[3][18] ), .S0(n860), .S1(n849), .Q(
        n790) );
  MUX41X1 U1065 ( .IN1(n790), .IN3(n788), .IN2(n789), .IN4(n787), .S0(n869), 
        .S1(n866), .Q(N38) );
  MUX41X1 U1066 ( .IN1(\regfile[12][19] ), .IN3(\regfile[14][19] ), .IN2(
        \regfile[13][19] ), .IN4(\regfile[15][19] ), .S0(n860), .S1(n849), .Q(
        n791) );
  MUX41X1 U1067 ( .IN1(\regfile[8][19] ), .IN3(\regfile[10][19] ), .IN2(
        \regfile[9][19] ), .IN4(\regfile[11][19] ), .S0(n860), .S1(n849), .Q(
        n792) );
  MUX41X1 U1068 ( .IN1(\regfile[4][19] ), .IN3(\regfile[6][19] ), .IN2(
        \regfile[5][19] ), .IN4(\regfile[7][19] ), .S0(n860), .S1(n849), .Q(
        n793) );
  MUX41X1 U1069 ( .IN1(\regfile[0][19] ), .IN3(\regfile[2][19] ), .IN2(
        \regfile[1][19] ), .IN4(\regfile[3][19] ), .S0(n860), .S1(n849), .Q(
        n794) );
  MUX41X1 U1070 ( .IN1(n794), .IN3(n792), .IN2(n793), .IN4(n791), .S0(n869), 
        .S1(n866), .Q(N37) );
  MUX41X1 U1071 ( .IN1(\regfile[12][20] ), .IN3(\regfile[14][20] ), .IN2(
        \regfile[13][20] ), .IN4(\regfile[15][20] ), .S0(n861), .S1(n850), .Q(
        n795) );
  MUX41X1 U1072 ( .IN1(\regfile[8][20] ), .IN3(\regfile[10][20] ), .IN2(
        \regfile[9][20] ), .IN4(\regfile[11][20] ), .S0(n861), .S1(n850), .Q(
        n796) );
  MUX41X1 U1073 ( .IN1(\regfile[4][20] ), .IN3(\regfile[6][20] ), .IN2(
        \regfile[5][20] ), .IN4(\regfile[7][20] ), .S0(n861), .S1(n850), .Q(
        n797) );
  MUX41X1 U1074 ( .IN1(\regfile[0][20] ), .IN3(\regfile[2][20] ), .IN2(
        \regfile[1][20] ), .IN4(\regfile[3][20] ), .S0(n861), .S1(n850), .Q(
        n798) );
  MUX41X1 U1075 ( .IN1(n798), .IN3(n796), .IN2(n797), .IN4(n795), .S0(n870), 
        .S1(n867), .Q(N36) );
  MUX41X1 U1076 ( .IN1(\regfile[12][21] ), .IN3(\regfile[14][21] ), .IN2(
        \regfile[13][21] ), .IN4(\regfile[15][21] ), .S0(n861), .S1(n850), .Q(
        n799) );
  MUX41X1 U1077 ( .IN1(\regfile[8][21] ), .IN3(\regfile[10][21] ), .IN2(
        \regfile[9][21] ), .IN4(\regfile[11][21] ), .S0(n861), .S1(n850), .Q(
        n800) );
  MUX41X1 U1078 ( .IN1(\regfile[4][21] ), .IN3(\regfile[6][21] ), .IN2(
        \regfile[5][21] ), .IN4(\regfile[7][21] ), .S0(n861), .S1(n850), .Q(
        n801) );
  MUX41X1 U1079 ( .IN1(\regfile[0][21] ), .IN3(\regfile[2][21] ), .IN2(
        \regfile[1][21] ), .IN4(\regfile[3][21] ), .S0(n861), .S1(n850), .Q(
        n802) );
  MUX41X1 U1080 ( .IN1(n802), .IN3(n800), .IN2(n801), .IN4(n799), .S0(n870), 
        .S1(n867), .Q(N35) );
  MUX41X1 U1081 ( .IN1(\regfile[12][22] ), .IN3(\regfile[14][22] ), .IN2(
        \regfile[13][22] ), .IN4(\regfile[15][22] ), .S0(n861), .S1(n850), .Q(
        n803) );
  MUX41X1 U1082 ( .IN1(\regfile[8][22] ), .IN3(\regfile[10][22] ), .IN2(
        \regfile[9][22] ), .IN4(\regfile[11][22] ), .S0(n861), .S1(n850), .Q(
        n804) );
  MUX41X1 U1083 ( .IN1(\regfile[4][22] ), .IN3(\regfile[6][22] ), .IN2(
        \regfile[5][22] ), .IN4(\regfile[7][22] ), .S0(n861), .S1(n850), .Q(
        n805) );
  MUX41X1 U1084 ( .IN1(\regfile[0][22] ), .IN3(\regfile[2][22] ), .IN2(
        \regfile[1][22] ), .IN4(\regfile[3][22] ), .S0(n861), .S1(n850), .Q(
        n806) );
  MUX41X1 U1085 ( .IN1(n806), .IN3(n804), .IN2(n805), .IN4(n803), .S0(n870), 
        .S1(n867), .Q(N34) );
  MUX41X1 U1086 ( .IN1(\regfile[12][23] ), .IN3(\regfile[14][23] ), .IN2(
        \regfile[13][23] ), .IN4(\regfile[15][23] ), .S0(n862), .S1(n851), .Q(
        n807) );
  MUX41X1 U1087 ( .IN1(\regfile[8][23] ), .IN3(\regfile[10][23] ), .IN2(
        \regfile[9][23] ), .IN4(\regfile[11][23] ), .S0(n862), .S1(n851), .Q(
        n808) );
  MUX41X1 U1088 ( .IN1(\regfile[4][23] ), .IN3(\regfile[6][23] ), .IN2(
        \regfile[5][23] ), .IN4(\regfile[7][23] ), .S0(n862), .S1(n851), .Q(
        n809) );
  MUX41X1 U1089 ( .IN1(\regfile[0][23] ), .IN3(\regfile[2][23] ), .IN2(
        \regfile[1][23] ), .IN4(\regfile[3][23] ), .S0(n862), .S1(n851), .Q(
        n810) );
  MUX41X1 U1090 ( .IN1(n810), .IN3(n808), .IN2(n809), .IN4(n807), .S0(n870), 
        .S1(n867), .Q(N33) );
  MUX41X1 U1091 ( .IN1(\regfile[12][24] ), .IN3(\regfile[14][24] ), .IN2(
        \regfile[13][24] ), .IN4(\regfile[15][24] ), .S0(n862), .S1(n851), .Q(
        n811) );
  MUX41X1 U1092 ( .IN1(\regfile[8][24] ), .IN3(\regfile[10][24] ), .IN2(
        \regfile[9][24] ), .IN4(\regfile[11][24] ), .S0(n862), .S1(n851), .Q(
        n812) );
  MUX41X1 U1093 ( .IN1(\regfile[4][24] ), .IN3(\regfile[6][24] ), .IN2(
        \regfile[5][24] ), .IN4(\regfile[7][24] ), .S0(n862), .S1(n851), .Q(
        n813) );
  MUX41X1 U1094 ( .IN1(\regfile[0][24] ), .IN3(\regfile[2][24] ), .IN2(
        \regfile[1][24] ), .IN4(\regfile[3][24] ), .S0(n862), .S1(n851), .Q(
        n814) );
  MUX41X1 U1095 ( .IN1(n814), .IN3(n812), .IN2(n813), .IN4(n811), .S0(n870), 
        .S1(n867), .Q(N32) );
  MUX41X1 U1096 ( .IN1(\regfile[12][25] ), .IN3(\regfile[14][25] ), .IN2(
        \regfile[13][25] ), .IN4(\regfile[15][25] ), .S0(n862), .S1(n851), .Q(
        n815) );
  MUX41X1 U1097 ( .IN1(\regfile[8][25] ), .IN3(\regfile[10][25] ), .IN2(
        \regfile[9][25] ), .IN4(\regfile[11][25] ), .S0(n862), .S1(n851), .Q(
        n816) );
  MUX41X1 U1098 ( .IN1(\regfile[4][25] ), .IN3(\regfile[6][25] ), .IN2(
        \regfile[5][25] ), .IN4(\regfile[7][25] ), .S0(n862), .S1(n851), .Q(
        n817) );
  MUX41X1 U1099 ( .IN1(\regfile[0][25] ), .IN3(\regfile[2][25] ), .IN2(
        \regfile[1][25] ), .IN4(\regfile[3][25] ), .S0(n862), .S1(n851), .Q(
        n818) );
  MUX41X1 U1100 ( .IN1(n818), .IN3(n816), .IN2(n817), .IN4(n815), .S0(n870), 
        .S1(n867), .Q(N31) );
  MUX41X1 U1101 ( .IN1(\regfile[12][26] ), .IN3(\regfile[14][26] ), .IN2(
        \regfile[13][26] ), .IN4(\regfile[15][26] ), .S0(n863), .S1(n852), .Q(
        n819) );
  MUX41X1 U1102 ( .IN1(\regfile[8][26] ), .IN3(\regfile[10][26] ), .IN2(
        \regfile[9][26] ), .IN4(\regfile[11][26] ), .S0(n863), .S1(n852), .Q(
        n820) );
  MUX41X1 U1103 ( .IN1(\regfile[4][26] ), .IN3(\regfile[6][26] ), .IN2(
        \regfile[5][26] ), .IN4(\regfile[7][26] ), .S0(n863), .S1(n852), .Q(
        n821) );
  MUX41X1 U1104 ( .IN1(\regfile[0][26] ), .IN3(\regfile[2][26] ), .IN2(
        \regfile[1][26] ), .IN4(\regfile[3][26] ), .S0(n863), .S1(n852), .Q(
        n822) );
  MUX41X1 U1105 ( .IN1(n822), .IN3(n820), .IN2(n821), .IN4(n819), .S0(n870), 
        .S1(n867), .Q(N30) );
  MUX41X1 U1106 ( .IN1(\regfile[12][27] ), .IN3(\regfile[14][27] ), .IN2(
        \regfile[13][27] ), .IN4(\regfile[15][27] ), .S0(n863), .S1(n852), .Q(
        n823) );
  MUX41X1 U1107 ( .IN1(\regfile[8][27] ), .IN3(\regfile[10][27] ), .IN2(
        \regfile[9][27] ), .IN4(\regfile[11][27] ), .S0(n863), .S1(n852), .Q(
        n824) );
  MUX41X1 U1108 ( .IN1(\regfile[4][27] ), .IN3(\regfile[6][27] ), .IN2(
        \regfile[5][27] ), .IN4(\regfile[7][27] ), .S0(n863), .S1(n852), .Q(
        n825) );
  MUX41X1 U1109 ( .IN1(\regfile[0][27] ), .IN3(\regfile[2][27] ), .IN2(
        \regfile[1][27] ), .IN4(\regfile[3][27] ), .S0(n863), .S1(n852), .Q(
        n826) );
  MUX41X1 U1110 ( .IN1(n826), .IN3(n824), .IN2(n825), .IN4(n823), .S0(n870), 
        .S1(n867), .Q(N29) );
  MUX41X1 U1111 ( .IN1(\regfile[12][28] ), .IN3(\regfile[14][28] ), .IN2(
        \regfile[13][28] ), .IN4(\regfile[15][28] ), .S0(n863), .S1(n852), .Q(
        n827) );
  MUX41X1 U1112 ( .IN1(\regfile[8][28] ), .IN3(\regfile[10][28] ), .IN2(
        \regfile[9][28] ), .IN4(\regfile[11][28] ), .S0(n863), .S1(n852), .Q(
        n828) );
  MUX41X1 U1113 ( .IN1(\regfile[4][28] ), .IN3(\regfile[6][28] ), .IN2(
        \regfile[5][28] ), .IN4(\regfile[7][28] ), .S0(n863), .S1(n852), .Q(
        n829) );
  MUX41X1 U1114 ( .IN1(\regfile[0][28] ), .IN3(\regfile[2][28] ), .IN2(
        \regfile[1][28] ), .IN4(\regfile[3][28] ), .S0(n863), .S1(n852), .Q(
        n830) );
  MUX41X1 U1115 ( .IN1(n830), .IN3(n828), .IN2(n829), .IN4(n827), .S0(n870), 
        .S1(n867), .Q(N28) );
  MUX41X1 U1116 ( .IN1(\regfile[12][29] ), .IN3(\regfile[14][29] ), .IN2(
        \regfile[13][29] ), .IN4(\regfile[15][29] ), .S0(n864), .S1(n853), .Q(
        n831) );
  MUX41X1 U1117 ( .IN1(\regfile[8][29] ), .IN3(\regfile[10][29] ), .IN2(
        \regfile[9][29] ), .IN4(\regfile[11][29] ), .S0(n864), .S1(n853), .Q(
        n832) );
  MUX41X1 U1118 ( .IN1(\regfile[4][29] ), .IN3(\regfile[6][29] ), .IN2(
        \regfile[5][29] ), .IN4(\regfile[7][29] ), .S0(n864), .S1(n853), .Q(
        n833) );
  MUX41X1 U1119 ( .IN1(\regfile[0][29] ), .IN3(\regfile[2][29] ), .IN2(
        \regfile[1][29] ), .IN4(\regfile[3][29] ), .S0(n864), .S1(n853), .Q(
        n834) );
  MUX41X1 U1120 ( .IN1(n834), .IN3(n832), .IN2(n833), .IN4(n831), .S0(n870), 
        .S1(n867), .Q(N27) );
  MUX41X1 U1121 ( .IN1(\regfile[12][30] ), .IN3(\regfile[14][30] ), .IN2(
        \regfile[13][30] ), .IN4(\regfile[15][30] ), .S0(n864), .S1(n853), .Q(
        n835) );
  MUX41X1 U1122 ( .IN1(\regfile[8][30] ), .IN3(\regfile[10][30] ), .IN2(
        \regfile[9][30] ), .IN4(\regfile[11][30] ), .S0(n864), .S1(n853), .Q(
        n836) );
  MUX41X1 U1123 ( .IN1(\regfile[4][30] ), .IN3(\regfile[6][30] ), .IN2(
        \regfile[5][30] ), .IN4(\regfile[7][30] ), .S0(n864), .S1(n853), .Q(
        n837) );
  MUX41X1 U1124 ( .IN1(\regfile[0][30] ), .IN3(\regfile[2][30] ), .IN2(
        \regfile[1][30] ), .IN4(\regfile[3][30] ), .S0(n864), .S1(n853), .Q(
        n838) );
  MUX41X1 U1125 ( .IN1(n838), .IN3(n836), .IN2(n837), .IN4(n835), .S0(n870), 
        .S1(n867), .Q(N26) );
  MUX41X1 U1126 ( .IN1(\regfile[12][31] ), .IN3(\regfile[14][31] ), .IN2(
        \regfile[13][31] ), .IN4(\regfile[15][31] ), .S0(n864), .S1(n853), .Q(
        n839) );
  MUX41X1 U1127 ( .IN1(\regfile[8][31] ), .IN3(\regfile[10][31] ), .IN2(
        \regfile[9][31] ), .IN4(\regfile[11][31] ), .S0(n864), .S1(n853), .Q(
        n840) );
  MUX41X1 U1128 ( .IN1(\regfile[4][31] ), .IN3(\regfile[6][31] ), .IN2(
        \regfile[5][31] ), .IN4(\regfile[7][31] ), .S0(n864), .S1(n853), .Q(
        n841) );
  MUX41X1 U1129 ( .IN1(\regfile[0][31] ), .IN3(\regfile[2][31] ), .IN2(
        \regfile[1][31] ), .IN4(\regfile[3][31] ), .S0(n864), .S1(n853), .Q(
        n842) );
  MUX41X1 U1130 ( .IN1(n842), .IN3(n840), .IN2(n841), .IN4(n839), .S0(n870), 
        .S1(n867), .Q(N25) );
  NBUFFX2 U1131 ( .INP(N18), .Z(n855) );
  NBUFFX2 U1132 ( .INP(N18), .Z(n856) );
  NBUFFX2 U1133 ( .INP(N18), .Z(n857) );
  NBUFFX2 U1134 ( .INP(N18), .Z(n858) );
  NBUFFX2 U1135 ( .INP(N18), .Z(n859) );
  NBUFFX2 U1136 ( .INP(N18), .Z(n860) );
  NBUFFX2 U1137 ( .INP(N18), .Z(n861) );
  NBUFFX2 U1138 ( .INP(N18), .Z(n862) );
  NBUFFX2 U1139 ( .INP(N18), .Z(n863) );
  NBUFFX2 U1140 ( .INP(N18), .Z(n864) );
  NBUFFX2 U1141 ( .INP(N20), .Z(n869) );
  NBUFFX2 U1142 ( .INP(N20), .Z(n870) );
  MUX41X1 U1143 ( .IN1(\regfile[12][0] ), .IN3(\regfile[14][0] ), .IN2(
        \regfile[13][0] ), .IN4(\regfile[15][0] ), .S0(n1010), .S1(n999), .Q(
        n871) );
  MUX41X1 U1144 ( .IN1(\regfile[8][0] ), .IN3(\regfile[10][0] ), .IN2(
        \regfile[9][0] ), .IN4(\regfile[11][0] ), .S0(n1010), .S1(n999), .Q(
        n872) );
  MUX41X1 U1145 ( .IN1(\regfile[4][0] ), .IN3(\regfile[6][0] ), .IN2(
        \regfile[5][0] ), .IN4(\regfile[7][0] ), .S0(n1010), .S1(n999), .Q(
        n873) );
  MUX41X1 U1146 ( .IN1(\regfile[0][0] ), .IN3(\regfile[2][0] ), .IN2(
        \regfile[1][0] ), .IN4(\regfile[3][0] ), .S0(n1010), .S1(n999), .Q(
        n874) );
  MUX41X1 U1147 ( .IN1(n874), .IN3(n872), .IN2(n873), .IN4(n871), .S0(n1024), 
        .S1(n1021), .Q(N88) );
  MUX41X1 U1148 ( .IN1(\regfile[12][1] ), .IN3(\regfile[14][1] ), .IN2(
        \regfile[13][1] ), .IN4(\regfile[15][1] ), .S0(n1010), .S1(n999), .Q(
        n875) );
  MUX41X1 U1149 ( .IN1(\regfile[8][1] ), .IN3(\regfile[10][1] ), .IN2(
        \regfile[9][1] ), .IN4(\regfile[11][1] ), .S0(n1010), .S1(n999), .Q(
        n876) );
  MUX41X1 U1150 ( .IN1(\regfile[4][1] ), .IN3(\regfile[6][1] ), .IN2(
        \regfile[5][1] ), .IN4(\regfile[7][1] ), .S0(n1010), .S1(n999), .Q(
        n877) );
  MUX41X1 U1151 ( .IN1(\regfile[0][1] ), .IN3(\regfile[2][1] ), .IN2(
        \regfile[1][1] ), .IN4(\regfile[3][1] ), .S0(n1010), .S1(n999), .Q(
        n878) );
  MUX41X1 U1152 ( .IN1(n878), .IN3(n876), .IN2(n877), .IN4(n875), .S0(n1024), 
        .S1(n1021), .Q(N87) );
  MUX41X1 U1153 ( .IN1(\regfile[12][2] ), .IN3(\regfile[14][2] ), .IN2(
        \regfile[13][2] ), .IN4(\regfile[15][2] ), .S0(n1011), .S1(n1000), .Q(
        n879) );
  MUX41X1 U1154 ( .IN1(\regfile[8][2] ), .IN3(\regfile[10][2] ), .IN2(
        \regfile[9][2] ), .IN4(\regfile[11][2] ), .S0(n1011), .S1(n1000), .Q(
        n880) );
  MUX41X1 U1155 ( .IN1(\regfile[4][2] ), .IN3(\regfile[6][2] ), .IN2(
        \regfile[5][2] ), .IN4(\regfile[7][2] ), .S0(n1011), .S1(n1000), .Q(
        n881) );
  MUX41X1 U1156 ( .IN1(\regfile[0][2] ), .IN3(\regfile[2][2] ), .IN2(
        \regfile[1][2] ), .IN4(\regfile[3][2] ), .S0(n1011), .S1(n1000), .Q(
        n882) );
  MUX41X1 U1157 ( .IN1(n882), .IN3(n880), .IN2(n881), .IN4(n879), .S0(n1024), 
        .S1(n1021), .Q(N86) );
  MUX41X1 U1158 ( .IN1(\regfile[12][3] ), .IN3(\regfile[14][3] ), .IN2(
        \regfile[13][3] ), .IN4(\regfile[15][3] ), .S0(n1011), .S1(n1000), .Q(
        n883) );
  MUX41X1 U1159 ( .IN1(\regfile[8][3] ), .IN3(\regfile[10][3] ), .IN2(
        \regfile[9][3] ), .IN4(\regfile[11][3] ), .S0(n1011), .S1(n1000), .Q(
        n884) );
  MUX41X1 U1160 ( .IN1(\regfile[4][3] ), .IN3(\regfile[6][3] ), .IN2(
        \regfile[5][3] ), .IN4(\regfile[7][3] ), .S0(n1011), .S1(n1000), .Q(
        n885) );
  MUX41X1 U1161 ( .IN1(\regfile[0][3] ), .IN3(\regfile[2][3] ), .IN2(
        \regfile[1][3] ), .IN4(\regfile[3][3] ), .S0(n1011), .S1(n1000), .Q(
        n886) );
  MUX41X1 U1162 ( .IN1(n886), .IN3(n884), .IN2(n885), .IN4(n883), .S0(n1024), 
        .S1(n1021), .Q(N85) );
  MUX41X1 U1163 ( .IN1(\regfile[12][4] ), .IN3(\regfile[14][4] ), .IN2(
        \regfile[13][4] ), .IN4(\regfile[15][4] ), .S0(n1011), .S1(n1000), .Q(
        n887) );
  MUX41X1 U1164 ( .IN1(\regfile[8][4] ), .IN3(\regfile[10][4] ), .IN2(
        \regfile[9][4] ), .IN4(\regfile[11][4] ), .S0(n1011), .S1(n1000), .Q(
        n888) );
  MUX41X1 U1165 ( .IN1(\regfile[4][4] ), .IN3(\regfile[6][4] ), .IN2(
        \regfile[5][4] ), .IN4(\regfile[7][4] ), .S0(n1011), .S1(n1000), .Q(
        n889) );
  MUX41X1 U1166 ( .IN1(\regfile[0][4] ), .IN3(\regfile[2][4] ), .IN2(
        \regfile[1][4] ), .IN4(\regfile[3][4] ), .S0(n1011), .S1(n1000), .Q(
        n890) );
  MUX41X1 U1167 ( .IN1(n890), .IN3(n888), .IN2(n889), .IN4(n887), .S0(n1024), 
        .S1(n1021), .Q(N84) );
  MUX41X1 U1168 ( .IN1(\regfile[12][5] ), .IN3(\regfile[14][5] ), .IN2(
        \regfile[13][5] ), .IN4(\regfile[15][5] ), .S0(n1012), .S1(n1001), .Q(
        n891) );
  MUX41X1 U1169 ( .IN1(\regfile[8][5] ), .IN3(\regfile[10][5] ), .IN2(
        \regfile[9][5] ), .IN4(\regfile[11][5] ), .S0(n1012), .S1(n1001), .Q(
        n892) );
  MUX41X1 U1170 ( .IN1(\regfile[4][5] ), .IN3(\regfile[6][5] ), .IN2(
        \regfile[5][5] ), .IN4(\regfile[7][5] ), .S0(n1012), .S1(n1001), .Q(
        n893) );
  MUX41X1 U1171 ( .IN1(\regfile[0][5] ), .IN3(\regfile[2][5] ), .IN2(
        \regfile[1][5] ), .IN4(\regfile[3][5] ), .S0(n1012), .S1(n1001), .Q(
        n894) );
  MUX41X1 U1172 ( .IN1(n894), .IN3(n892), .IN2(n893), .IN4(n891), .S0(n1024), 
        .S1(n1021), .Q(N83) );
  MUX41X1 U1173 ( .IN1(\regfile[12][6] ), .IN3(\regfile[14][6] ), .IN2(
        \regfile[13][6] ), .IN4(\regfile[15][6] ), .S0(n1012), .S1(n1001), .Q(
        n895) );
  MUX41X1 U1174 ( .IN1(\regfile[8][6] ), .IN3(\regfile[10][6] ), .IN2(
        \regfile[9][6] ), .IN4(\regfile[11][6] ), .S0(n1012), .S1(n1001), .Q(
        n896) );
  MUX41X1 U1175 ( .IN1(\regfile[4][6] ), .IN3(\regfile[6][6] ), .IN2(
        \regfile[5][6] ), .IN4(\regfile[7][6] ), .S0(n1012), .S1(n1001), .Q(
        n897) );
  MUX41X1 U1176 ( .IN1(\regfile[0][6] ), .IN3(\regfile[2][6] ), .IN2(
        \regfile[1][6] ), .IN4(\regfile[3][6] ), .S0(n1012), .S1(n1001), .Q(
        n898) );
  MUX41X1 U1177 ( .IN1(n898), .IN3(n896), .IN2(n897), .IN4(n895), .S0(n1024), 
        .S1(n1021), .Q(N82) );
  MUX41X1 U1178 ( .IN1(\regfile[12][7] ), .IN3(\regfile[14][7] ), .IN2(
        \regfile[13][7] ), .IN4(\regfile[15][7] ), .S0(n1012), .S1(n1001), .Q(
        n899) );
  MUX41X1 U1179 ( .IN1(\regfile[8][7] ), .IN3(\regfile[10][7] ), .IN2(
        \regfile[9][7] ), .IN4(\regfile[11][7] ), .S0(n1012), .S1(n1001), .Q(
        n900) );
  MUX41X1 U1180 ( .IN1(\regfile[4][7] ), .IN3(\regfile[6][7] ), .IN2(
        \regfile[5][7] ), .IN4(\regfile[7][7] ), .S0(n1012), .S1(n1001), .Q(
        n901) );
  MUX41X1 U1181 ( .IN1(\regfile[0][7] ), .IN3(\regfile[2][7] ), .IN2(
        \regfile[1][7] ), .IN4(\regfile[3][7] ), .S0(n1012), .S1(n1001), .Q(
        n902) );
  MUX41X1 U1182 ( .IN1(n902), .IN3(n900), .IN2(n901), .IN4(n899), .S0(n1024), 
        .S1(n1021), .Q(N81) );
  MUX41X1 U1183 ( .IN1(\regfile[12][8] ), .IN3(\regfile[14][8] ), .IN2(
        \regfile[13][8] ), .IN4(\regfile[15][8] ), .S0(n1013), .S1(n1002), .Q(
        n903) );
  MUX41X1 U1184 ( .IN1(\regfile[8][8] ), .IN3(\regfile[10][8] ), .IN2(
        \regfile[9][8] ), .IN4(\regfile[11][8] ), .S0(n1013), .S1(n1002), .Q(
        n904) );
  MUX41X1 U1185 ( .IN1(\regfile[4][8] ), .IN3(\regfile[6][8] ), .IN2(
        \regfile[5][8] ), .IN4(\regfile[7][8] ), .S0(n1013), .S1(n1002), .Q(
        n905) );
  MUX41X1 U1186 ( .IN1(\regfile[0][8] ), .IN3(\regfile[2][8] ), .IN2(
        \regfile[1][8] ), .IN4(\regfile[3][8] ), .S0(n1013), .S1(n1002), .Q(
        n906) );
  MUX41X1 U1187 ( .IN1(n906), .IN3(n904), .IN2(n905), .IN4(n903), .S0(n1025), 
        .S1(n1022), .Q(N80) );
  MUX41X1 U1188 ( .IN1(\regfile[12][9] ), .IN3(\regfile[14][9] ), .IN2(
        \regfile[13][9] ), .IN4(\regfile[15][9] ), .S0(n1013), .S1(n1002), .Q(
        n907) );
  MUX41X1 U1189 ( .IN1(\regfile[8][9] ), .IN3(\regfile[10][9] ), .IN2(
        \regfile[9][9] ), .IN4(\regfile[11][9] ), .S0(n1013), .S1(n1002), .Q(
        n908) );
  MUX41X1 U1190 ( .IN1(\regfile[4][9] ), .IN3(\regfile[6][9] ), .IN2(
        \regfile[5][9] ), .IN4(\regfile[7][9] ), .S0(n1013), .S1(n1002), .Q(
        n909) );
  MUX41X1 U1191 ( .IN1(\regfile[0][9] ), .IN3(\regfile[2][9] ), .IN2(
        \regfile[1][9] ), .IN4(\regfile[3][9] ), .S0(n1013), .S1(n1002), .Q(
        n910) );
  MUX41X1 U1192 ( .IN1(n910), .IN3(n908), .IN2(n909), .IN4(n907), .S0(n1025), 
        .S1(n1022), .Q(N79) );
  MUX41X1 U1193 ( .IN1(\regfile[12][10] ), .IN3(\regfile[14][10] ), .IN2(
        \regfile[13][10] ), .IN4(\regfile[15][10] ), .S0(n1013), .S1(n1002), 
        .Q(n911) );
  MUX41X1 U1194 ( .IN1(\regfile[8][10] ), .IN3(\regfile[10][10] ), .IN2(
        \regfile[9][10] ), .IN4(\regfile[11][10] ), .S0(n1013), .S1(n1002), 
        .Q(n912) );
  MUX41X1 U1195 ( .IN1(\regfile[4][10] ), .IN3(\regfile[6][10] ), .IN2(
        \regfile[5][10] ), .IN4(\regfile[7][10] ), .S0(n1013), .S1(n1002), .Q(
        n913) );
  MUX41X1 U1196 ( .IN1(\regfile[0][10] ), .IN3(\regfile[2][10] ), .IN2(
        \regfile[1][10] ), .IN4(\regfile[3][10] ), .S0(n1013), .S1(n1002), .Q(
        n914) );
  MUX41X1 U1197 ( .IN1(n914), .IN3(n912), .IN2(n913), .IN4(n911), .S0(n1025), 
        .S1(n1022), .Q(N78) );
  MUX41X1 U1198 ( .IN1(\regfile[12][11] ), .IN3(\regfile[14][11] ), .IN2(
        \regfile[13][11] ), .IN4(\regfile[15][11] ), .S0(n1014), .S1(n1003), 
        .Q(n915) );
  MUX41X1 U1199 ( .IN1(\regfile[8][11] ), .IN3(\regfile[10][11] ), .IN2(
        \regfile[9][11] ), .IN4(\regfile[11][11] ), .S0(n1014), .S1(n1003), 
        .Q(n916) );
  MUX41X1 U1200 ( .IN1(\regfile[4][11] ), .IN3(\regfile[6][11] ), .IN2(
        \regfile[5][11] ), .IN4(\regfile[7][11] ), .S0(n1014), .S1(n1003), .Q(
        n917) );
  MUX41X1 U1201 ( .IN1(\regfile[0][11] ), .IN3(\regfile[2][11] ), .IN2(
        \regfile[1][11] ), .IN4(\regfile[3][11] ), .S0(n1014), .S1(n1003), .Q(
        n918) );
  MUX41X1 U1202 ( .IN1(n918), .IN3(n916), .IN2(n917), .IN4(n915), .S0(n1025), 
        .S1(n1022), .Q(N77) );
  MUX41X1 U1203 ( .IN1(\regfile[12][12] ), .IN3(\regfile[14][12] ), .IN2(
        \regfile[13][12] ), .IN4(\regfile[15][12] ), .S0(n1014), .S1(n1003), 
        .Q(n919) );
  MUX41X1 U1204 ( .IN1(\regfile[8][12] ), .IN3(\regfile[10][12] ), .IN2(
        \regfile[9][12] ), .IN4(\regfile[11][12] ), .S0(n1014), .S1(n1003), 
        .Q(n920) );
  MUX41X1 U1205 ( .IN1(\regfile[4][12] ), .IN3(\regfile[6][12] ), .IN2(
        \regfile[5][12] ), .IN4(\regfile[7][12] ), .S0(n1014), .S1(n1003), .Q(
        n921) );
  MUX41X1 U1206 ( .IN1(\regfile[0][12] ), .IN3(\regfile[2][12] ), .IN2(
        \regfile[1][12] ), .IN4(\regfile[3][12] ), .S0(n1014), .S1(n1003), .Q(
        n922) );
  MUX41X1 U1207 ( .IN1(n922), .IN3(n920), .IN2(n921), .IN4(n919), .S0(n1025), 
        .S1(n1022), .Q(N76) );
  MUX41X1 U1208 ( .IN1(\regfile[12][13] ), .IN3(\regfile[14][13] ), .IN2(
        \regfile[13][13] ), .IN4(\regfile[15][13] ), .S0(n1014), .S1(n1003), 
        .Q(n923) );
  MUX41X1 U1209 ( .IN1(\regfile[8][13] ), .IN3(\regfile[10][13] ), .IN2(
        \regfile[9][13] ), .IN4(\regfile[11][13] ), .S0(n1014), .S1(n1003), 
        .Q(n924) );
  MUX41X1 U1210 ( .IN1(\regfile[4][13] ), .IN3(\regfile[6][13] ), .IN2(
        \regfile[5][13] ), .IN4(\regfile[7][13] ), .S0(n1014), .S1(n1003), .Q(
        n925) );
  MUX41X1 U1211 ( .IN1(\regfile[0][13] ), .IN3(\regfile[2][13] ), .IN2(
        \regfile[1][13] ), .IN4(\regfile[3][13] ), .S0(n1014), .S1(n1003), .Q(
        n926) );
  MUX41X1 U1212 ( .IN1(n926), .IN3(n924), .IN2(n925), .IN4(n923), .S0(n1025), 
        .S1(n1022), .Q(N75) );
  MUX41X1 U1213 ( .IN1(\regfile[12][14] ), .IN3(\regfile[14][14] ), .IN2(
        \regfile[13][14] ), .IN4(\regfile[15][14] ), .S0(n1015), .S1(n1004), 
        .Q(n927) );
  MUX41X1 U1214 ( .IN1(\regfile[8][14] ), .IN3(\regfile[10][14] ), .IN2(
        \regfile[9][14] ), .IN4(\regfile[11][14] ), .S0(n1015), .S1(n1004), 
        .Q(n928) );
  MUX41X1 U1215 ( .IN1(\regfile[4][14] ), .IN3(\regfile[6][14] ), .IN2(
        \regfile[5][14] ), .IN4(\regfile[7][14] ), .S0(n1015), .S1(n1004), .Q(
        n929) );
  MUX41X1 U1216 ( .IN1(\regfile[0][14] ), .IN3(\regfile[2][14] ), .IN2(
        \regfile[1][14] ), .IN4(\regfile[3][14] ), .S0(n1015), .S1(n1004), .Q(
        n930) );
  MUX41X1 U1217 ( .IN1(n930), .IN3(n928), .IN2(n929), .IN4(n927), .S0(n1025), 
        .S1(n1022), .Q(N74) );
  MUX41X1 U1218 ( .IN1(\regfile[12][15] ), .IN3(\regfile[14][15] ), .IN2(
        \regfile[13][15] ), .IN4(\regfile[15][15] ), .S0(n1015), .S1(n1004), 
        .Q(n931) );
  MUX41X1 U1219 ( .IN1(\regfile[8][15] ), .IN3(\regfile[10][15] ), .IN2(
        \regfile[9][15] ), .IN4(\regfile[11][15] ), .S0(n1015), .S1(n1004), 
        .Q(n932) );
  MUX41X1 U1220 ( .IN1(\regfile[4][15] ), .IN3(\regfile[6][15] ), .IN2(
        \regfile[5][15] ), .IN4(\regfile[7][15] ), .S0(n1015), .S1(n1004), .Q(
        n933) );
  MUX41X1 U1221 ( .IN1(\regfile[0][15] ), .IN3(\regfile[2][15] ), .IN2(
        \regfile[1][15] ), .IN4(\regfile[3][15] ), .S0(n1015), .S1(n1004), .Q(
        n934) );
  MUX41X1 U1222 ( .IN1(n934), .IN3(n932), .IN2(n933), .IN4(n931), .S0(n1025), 
        .S1(n1022), .Q(N73) );
  MUX41X1 U1223 ( .IN1(\regfile[12][16] ), .IN3(\regfile[14][16] ), .IN2(
        \regfile[13][16] ), .IN4(\regfile[15][16] ), .S0(n1015), .S1(n1004), 
        .Q(n935) );
  MUX41X1 U1224 ( .IN1(\regfile[8][16] ), .IN3(\regfile[10][16] ), .IN2(
        \regfile[9][16] ), .IN4(\regfile[11][16] ), .S0(n1015), .S1(n1004), 
        .Q(n936) );
  MUX41X1 U1225 ( .IN1(\regfile[4][16] ), .IN3(\regfile[6][16] ), .IN2(
        \regfile[5][16] ), .IN4(\regfile[7][16] ), .S0(n1015), .S1(n1004), .Q(
        n937) );
  MUX41X1 U1226 ( .IN1(\regfile[0][16] ), .IN3(\regfile[2][16] ), .IN2(
        \regfile[1][16] ), .IN4(\regfile[3][16] ), .S0(n1015), .S1(n1004), .Q(
        n938) );
  MUX41X1 U1227 ( .IN1(n938), .IN3(n936), .IN2(n937), .IN4(n935), .S0(n1025), 
        .S1(n1022), .Q(N72) );
  MUX41X1 U1228 ( .IN1(\regfile[12][17] ), .IN3(\regfile[14][17] ), .IN2(
        \regfile[13][17] ), .IN4(\regfile[15][17] ), .S0(n1016), .S1(n1005), 
        .Q(n939) );
  MUX41X1 U1229 ( .IN1(\regfile[8][17] ), .IN3(\regfile[10][17] ), .IN2(
        \regfile[9][17] ), .IN4(\regfile[11][17] ), .S0(n1016), .S1(n1005), 
        .Q(n940) );
  MUX41X1 U1230 ( .IN1(\regfile[4][17] ), .IN3(\regfile[6][17] ), .IN2(
        \regfile[5][17] ), .IN4(\regfile[7][17] ), .S0(n1016), .S1(n1005), .Q(
        n941) );
  MUX41X1 U1231 ( .IN1(\regfile[0][17] ), .IN3(\regfile[2][17] ), .IN2(
        \regfile[1][17] ), .IN4(\regfile[3][17] ), .S0(n1016), .S1(n1005), .Q(
        n942) );
  MUX41X1 U1232 ( .IN1(n942), .IN3(n940), .IN2(n941), .IN4(n939), .S0(n1025), 
        .S1(n1022), .Q(N71) );
  MUX41X1 U1233 ( .IN1(\regfile[12][18] ), .IN3(\regfile[14][18] ), .IN2(
        \regfile[13][18] ), .IN4(\regfile[15][18] ), .S0(n1016), .S1(n1005), 
        .Q(n943) );
  MUX41X1 U1234 ( .IN1(\regfile[8][18] ), .IN3(\regfile[10][18] ), .IN2(
        \regfile[9][18] ), .IN4(\regfile[11][18] ), .S0(n1016), .S1(n1005), 
        .Q(n944) );
  MUX41X1 U1235 ( .IN1(\regfile[4][18] ), .IN3(\regfile[6][18] ), .IN2(
        \regfile[5][18] ), .IN4(\regfile[7][18] ), .S0(n1016), .S1(n1005), .Q(
        n945) );
  MUX41X1 U1236 ( .IN1(\regfile[0][18] ), .IN3(\regfile[2][18] ), .IN2(
        \regfile[1][18] ), .IN4(\regfile[3][18] ), .S0(n1016), .S1(n1005), .Q(
        n946) );
  MUX41X1 U1237 ( .IN1(n946), .IN3(n944), .IN2(n945), .IN4(n943), .S0(n1025), 
        .S1(n1022), .Q(N70) );
  MUX41X1 U1238 ( .IN1(\regfile[12][19] ), .IN3(\regfile[14][19] ), .IN2(
        \regfile[13][19] ), .IN4(\regfile[15][19] ), .S0(n1016), .S1(n1005), 
        .Q(n947) );
  MUX41X1 U1239 ( .IN1(\regfile[8][19] ), .IN3(\regfile[10][19] ), .IN2(
        \regfile[9][19] ), .IN4(\regfile[11][19] ), .S0(n1016), .S1(n1005), 
        .Q(n948) );
  MUX41X1 U1240 ( .IN1(\regfile[4][19] ), .IN3(\regfile[6][19] ), .IN2(
        \regfile[5][19] ), .IN4(\regfile[7][19] ), .S0(n1016), .S1(n1005), .Q(
        n949) );
  MUX41X1 U1241 ( .IN1(\regfile[0][19] ), .IN3(\regfile[2][19] ), .IN2(
        \regfile[1][19] ), .IN4(\regfile[3][19] ), .S0(n1016), .S1(n1005), .Q(
        n950) );
  MUX41X1 U1242 ( .IN1(n950), .IN3(n948), .IN2(n949), .IN4(n947), .S0(n1025), 
        .S1(n1022), .Q(N69) );
  MUX41X1 U1243 ( .IN1(\regfile[12][20] ), .IN3(\regfile[14][20] ), .IN2(
        \regfile[13][20] ), .IN4(\regfile[15][20] ), .S0(n1017), .S1(n1006), 
        .Q(n951) );
  MUX41X1 U1244 ( .IN1(\regfile[8][20] ), .IN3(\regfile[10][20] ), .IN2(
        \regfile[9][20] ), .IN4(\regfile[11][20] ), .S0(n1017), .S1(n1006), 
        .Q(n952) );
  MUX41X1 U1245 ( .IN1(\regfile[4][20] ), .IN3(\regfile[6][20] ), .IN2(
        \regfile[5][20] ), .IN4(\regfile[7][20] ), .S0(n1017), .S1(n1006), .Q(
        n953) );
  MUX41X1 U1246 ( .IN1(\regfile[0][20] ), .IN3(\regfile[2][20] ), .IN2(
        \regfile[1][20] ), .IN4(\regfile[3][20] ), .S0(n1017), .S1(n1006), .Q(
        n954) );
  MUX41X1 U1247 ( .IN1(n954), .IN3(n952), .IN2(n953), .IN4(n951), .S0(n1026), 
        .S1(n1023), .Q(N68) );
  MUX41X1 U1248 ( .IN1(\regfile[12][21] ), .IN3(\regfile[14][21] ), .IN2(
        \regfile[13][21] ), .IN4(\regfile[15][21] ), .S0(n1017), .S1(n1006), 
        .Q(n955) );
  MUX41X1 U1249 ( .IN1(\regfile[8][21] ), .IN3(\regfile[10][21] ), .IN2(
        \regfile[9][21] ), .IN4(\regfile[11][21] ), .S0(n1017), .S1(n1006), 
        .Q(n956) );
  MUX41X1 U1250 ( .IN1(\regfile[4][21] ), .IN3(\regfile[6][21] ), .IN2(
        \regfile[5][21] ), .IN4(\regfile[7][21] ), .S0(n1017), .S1(n1006), .Q(
        n957) );
  MUX41X1 U1251 ( .IN1(\regfile[0][21] ), .IN3(\regfile[2][21] ), .IN2(
        \regfile[1][21] ), .IN4(\regfile[3][21] ), .S0(n1017), .S1(n1006), .Q(
        n958) );
  MUX41X1 U1252 ( .IN1(n958), .IN3(n956), .IN2(n957), .IN4(n955), .S0(n1026), 
        .S1(n1023), .Q(N67) );
  MUX41X1 U1253 ( .IN1(\regfile[12][22] ), .IN3(\regfile[14][22] ), .IN2(
        \regfile[13][22] ), .IN4(\regfile[15][22] ), .S0(n1017), .S1(n1006), 
        .Q(n959) );
  MUX41X1 U1254 ( .IN1(\regfile[8][22] ), .IN3(\regfile[10][22] ), .IN2(
        \regfile[9][22] ), .IN4(\regfile[11][22] ), .S0(n1017), .S1(n1006), 
        .Q(n960) );
  MUX41X1 U1255 ( .IN1(\regfile[4][22] ), .IN3(\regfile[6][22] ), .IN2(
        \regfile[5][22] ), .IN4(\regfile[7][22] ), .S0(n1017), .S1(n1006), .Q(
        n961) );
  MUX41X1 U1256 ( .IN1(\regfile[0][22] ), .IN3(\regfile[2][22] ), .IN2(
        \regfile[1][22] ), .IN4(\regfile[3][22] ), .S0(n1017), .S1(n1006), .Q(
        n962) );
  MUX41X1 U1257 ( .IN1(n962), .IN3(n960), .IN2(n961), .IN4(n959), .S0(n1026), 
        .S1(n1023), .Q(N66) );
  MUX41X1 U1258 ( .IN1(\regfile[12][23] ), .IN3(\regfile[14][23] ), .IN2(
        \regfile[13][23] ), .IN4(\regfile[15][23] ), .S0(n1018), .S1(n1007), 
        .Q(n963) );
  MUX41X1 U1259 ( .IN1(\regfile[8][23] ), .IN3(\regfile[10][23] ), .IN2(
        \regfile[9][23] ), .IN4(\regfile[11][23] ), .S0(n1018), .S1(n1007), 
        .Q(n964) );
  MUX41X1 U1260 ( .IN1(\regfile[4][23] ), .IN3(\regfile[6][23] ), .IN2(
        \regfile[5][23] ), .IN4(\regfile[7][23] ), .S0(n1018), .S1(n1007), .Q(
        n965) );
  MUX41X1 U1261 ( .IN1(\regfile[0][23] ), .IN3(\regfile[2][23] ), .IN2(
        \regfile[1][23] ), .IN4(\regfile[3][23] ), .S0(n1018), .S1(n1007), .Q(
        n966) );
  MUX41X1 U1262 ( .IN1(n966), .IN3(n964), .IN2(n965), .IN4(n963), .S0(n1026), 
        .S1(n1023), .Q(N65) );
  MUX41X1 U1263 ( .IN1(\regfile[12][24] ), .IN3(\regfile[14][24] ), .IN2(
        \regfile[13][24] ), .IN4(\regfile[15][24] ), .S0(n1018), .S1(n1007), 
        .Q(n967) );
  MUX41X1 U1264 ( .IN1(\regfile[8][24] ), .IN3(\regfile[10][24] ), .IN2(
        \regfile[9][24] ), .IN4(\regfile[11][24] ), .S0(n1018), .S1(n1007), 
        .Q(n968) );
  MUX41X1 U1265 ( .IN1(\regfile[4][24] ), .IN3(\regfile[6][24] ), .IN2(
        \regfile[5][24] ), .IN4(\regfile[7][24] ), .S0(n1018), .S1(n1007), .Q(
        n969) );
  MUX41X1 U1266 ( .IN1(\regfile[0][24] ), .IN3(\regfile[2][24] ), .IN2(
        \regfile[1][24] ), .IN4(\regfile[3][24] ), .S0(n1018), .S1(n1007), .Q(
        n970) );
  MUX41X1 U1267 ( .IN1(n970), .IN3(n968), .IN2(n969), .IN4(n967), .S0(n1026), 
        .S1(n1023), .Q(N64) );
  MUX41X1 U1268 ( .IN1(\regfile[12][25] ), .IN3(\regfile[14][25] ), .IN2(
        \regfile[13][25] ), .IN4(\regfile[15][25] ), .S0(n1018), .S1(n1007), 
        .Q(n971) );
  MUX41X1 U1269 ( .IN1(\regfile[8][25] ), .IN3(\regfile[10][25] ), .IN2(
        \regfile[9][25] ), .IN4(\regfile[11][25] ), .S0(n1018), .S1(n1007), 
        .Q(n972) );
  MUX41X1 U1270 ( .IN1(\regfile[4][25] ), .IN3(\regfile[6][25] ), .IN2(
        \regfile[5][25] ), .IN4(\regfile[7][25] ), .S0(n1018), .S1(n1007), .Q(
        n973) );
  MUX41X1 U1271 ( .IN1(\regfile[0][25] ), .IN3(\regfile[2][25] ), .IN2(
        \regfile[1][25] ), .IN4(\regfile[3][25] ), .S0(n1018), .S1(n1007), .Q(
        n974) );
  MUX41X1 U1272 ( .IN1(n974), .IN3(n972), .IN2(n973), .IN4(n971), .S0(n1026), 
        .S1(n1023), .Q(N63) );
  MUX41X1 U1273 ( .IN1(\regfile[12][26] ), .IN3(\regfile[14][26] ), .IN2(
        \regfile[13][26] ), .IN4(\regfile[15][26] ), .S0(n1019), .S1(n1008), 
        .Q(n975) );
  MUX41X1 U1274 ( .IN1(\regfile[8][26] ), .IN3(\regfile[10][26] ), .IN2(
        \regfile[9][26] ), .IN4(\regfile[11][26] ), .S0(n1019), .S1(n1008), 
        .Q(n976) );
  MUX41X1 U1275 ( .IN1(\regfile[4][26] ), .IN3(\regfile[6][26] ), .IN2(
        \regfile[5][26] ), .IN4(\regfile[7][26] ), .S0(n1019), .S1(n1008), .Q(
        n977) );
  MUX41X1 U1276 ( .IN1(\regfile[0][26] ), .IN3(\regfile[2][26] ), .IN2(
        \regfile[1][26] ), .IN4(\regfile[3][26] ), .S0(n1019), .S1(n1008), .Q(
        n978) );
  MUX41X1 U1277 ( .IN1(n978), .IN3(n976), .IN2(n977), .IN4(n975), .S0(n1026), 
        .S1(n1023), .Q(N62) );
  MUX41X1 U1278 ( .IN1(\regfile[12][27] ), .IN3(\regfile[14][27] ), .IN2(
        \regfile[13][27] ), .IN4(\regfile[15][27] ), .S0(n1019), .S1(n1008), 
        .Q(n979) );
  MUX41X1 U1279 ( .IN1(\regfile[8][27] ), .IN3(\regfile[10][27] ), .IN2(
        \regfile[9][27] ), .IN4(\regfile[11][27] ), .S0(n1019), .S1(n1008), 
        .Q(n980) );
  MUX41X1 U1280 ( .IN1(\regfile[4][27] ), .IN3(\regfile[6][27] ), .IN2(
        \regfile[5][27] ), .IN4(\regfile[7][27] ), .S0(n1019), .S1(n1008), .Q(
        n981) );
  MUX41X1 U1281 ( .IN1(\regfile[0][27] ), .IN3(\regfile[2][27] ), .IN2(
        \regfile[1][27] ), .IN4(\regfile[3][27] ), .S0(n1019), .S1(n1008), .Q(
        n982) );
  MUX41X1 U1282 ( .IN1(n982), .IN3(n980), .IN2(n981), .IN4(n979), .S0(n1026), 
        .S1(n1023), .Q(N61) );
  MUX41X1 U1283 ( .IN1(\regfile[12][28] ), .IN3(\regfile[14][28] ), .IN2(
        \regfile[13][28] ), .IN4(\regfile[15][28] ), .S0(n1019), .S1(n1008), 
        .Q(n983) );
  MUX41X1 U1284 ( .IN1(\regfile[8][28] ), .IN3(\regfile[10][28] ), .IN2(
        \regfile[9][28] ), .IN4(\regfile[11][28] ), .S0(n1019), .S1(n1008), 
        .Q(n984) );
  MUX41X1 U1285 ( .IN1(\regfile[4][28] ), .IN3(\regfile[6][28] ), .IN2(
        \regfile[5][28] ), .IN4(\regfile[7][28] ), .S0(n1019), .S1(n1008), .Q(
        n985) );
  MUX41X1 U1286 ( .IN1(\regfile[0][28] ), .IN3(\regfile[2][28] ), .IN2(
        \regfile[1][28] ), .IN4(\regfile[3][28] ), .S0(n1019), .S1(n1008), .Q(
        n986) );
  MUX41X1 U1287 ( .IN1(n986), .IN3(n984), .IN2(n985), .IN4(n983), .S0(n1026), 
        .S1(n1023), .Q(N60) );
  MUX41X1 U1288 ( .IN1(\regfile[12][29] ), .IN3(\regfile[14][29] ), .IN2(
        \regfile[13][29] ), .IN4(\regfile[15][29] ), .S0(n1020), .S1(n1009), 
        .Q(n987) );
  MUX41X1 U1289 ( .IN1(\regfile[8][29] ), .IN3(\regfile[10][29] ), .IN2(
        \regfile[9][29] ), .IN4(\regfile[11][29] ), .S0(n1020), .S1(n1009), 
        .Q(n988) );
  MUX41X1 U1290 ( .IN1(\regfile[4][29] ), .IN3(\regfile[6][29] ), .IN2(
        \regfile[5][29] ), .IN4(\regfile[7][29] ), .S0(n1020), .S1(n1009), .Q(
        n989) );
  MUX41X1 U1291 ( .IN1(\regfile[0][29] ), .IN3(\regfile[2][29] ), .IN2(
        \regfile[1][29] ), .IN4(\regfile[3][29] ), .S0(n1020), .S1(n1009), .Q(
        n990) );
  MUX41X1 U1292 ( .IN1(n990), .IN3(n988), .IN2(n989), .IN4(n987), .S0(n1026), 
        .S1(n1023), .Q(N59) );
  MUX41X1 U1293 ( .IN1(\regfile[12][30] ), .IN3(\regfile[14][30] ), .IN2(
        \regfile[13][30] ), .IN4(\regfile[15][30] ), .S0(n1020), .S1(n1009), 
        .Q(n991) );
  MUX41X1 U1294 ( .IN1(\regfile[8][30] ), .IN3(\regfile[10][30] ), .IN2(
        \regfile[9][30] ), .IN4(\regfile[11][30] ), .S0(n1020), .S1(n1009), 
        .Q(n992) );
  MUX41X1 U1295 ( .IN1(\regfile[4][30] ), .IN3(\regfile[6][30] ), .IN2(
        \regfile[5][30] ), .IN4(\regfile[7][30] ), .S0(n1020), .S1(n1009), .Q(
        n993) );
  MUX41X1 U1296 ( .IN1(\regfile[0][30] ), .IN3(\regfile[2][30] ), .IN2(
        \regfile[1][30] ), .IN4(\regfile[3][30] ), .S0(n1020), .S1(n1009), .Q(
        n994) );
  MUX41X1 U1297 ( .IN1(n994), .IN3(n992), .IN2(n993), .IN4(n991), .S0(n1026), 
        .S1(n1023), .Q(N58) );
  MUX41X1 U1298 ( .IN1(\regfile[12][31] ), .IN3(\regfile[14][31] ), .IN2(
        \regfile[13][31] ), .IN4(\regfile[15][31] ), .S0(n1020), .S1(n1009), 
        .Q(n995) );
  MUX41X1 U1299 ( .IN1(\regfile[8][31] ), .IN3(\regfile[10][31] ), .IN2(
        \regfile[9][31] ), .IN4(\regfile[11][31] ), .S0(n1020), .S1(n1009), 
        .Q(n996) );
  MUX41X1 U1300 ( .IN1(\regfile[4][31] ), .IN3(\regfile[6][31] ), .IN2(
        \regfile[5][31] ), .IN4(\regfile[7][31] ), .S0(n1020), .S1(n1009), .Q(
        n997) );
  MUX41X1 U1301 ( .IN1(\regfile[0][31] ), .IN3(\regfile[2][31] ), .IN2(
        \regfile[1][31] ), .IN4(\regfile[3][31] ), .S0(n1020), .S1(n1009), .Q(
        n998) );
  MUX41X1 U1302 ( .IN1(n998), .IN3(n996), .IN2(n997), .IN4(n995), .S0(n1026), 
        .S1(n1023), .Q(N57) );
  NBUFFX2 U1303 ( .INP(N22), .Z(n1011) );
  NBUFFX2 U1304 ( .INP(N22), .Z(n1012) );
  NBUFFX2 U1305 ( .INP(N22), .Z(n1013) );
  NBUFFX2 U1306 ( .INP(N22), .Z(n1014) );
  NBUFFX2 U1307 ( .INP(N22), .Z(n1015) );
  NBUFFX2 U1308 ( .INP(N22), .Z(n1016) );
  NBUFFX2 U1309 ( .INP(N22), .Z(n1017) );
  NBUFFX2 U1310 ( .INP(N22), .Z(n1018) );
  NBUFFX2 U1311 ( .INP(N22), .Z(n1019) );
  NBUFFX2 U1312 ( .INP(N22), .Z(n1020) );
  NBUFFX2 U1313 ( .INP(N24), .Z(n1025) );
  NBUFFX2 U1314 ( .INP(N24), .Z(n1026) );
  NBUFFX2 U1315 ( .INP(n1172), .Z(n1027) );
  NBUFFX2 U1316 ( .INP(n1172), .Z(n1028) );
  NBUFFX2 U1317 ( .INP(n1172), .Z(n1029) );
  NBUFFX2 U1318 ( .INP(n1172), .Z(n1030) );
  NBUFFX2 U1319 ( .INP(n1172), .Z(n1031) );
  NBUFFX2 U1320 ( .INP(n80), .Z(n1032) );
  NBUFFX2 U1321 ( .INP(n78), .Z(n1033) );
  NBUFFX2 U1322 ( .INP(n78), .Z(n1034) );
  NBUFFX2 U1323 ( .INP(n70), .Z(n1036) );
  NBUFFX2 U1324 ( .INP(n70), .Z(n1037) );
  NBUFFX2 U1325 ( .INP(n68), .Z(n1039) );
  NBUFFX2 U1326 ( .INP(n68), .Z(n1040) );
  INVX0 U1327 ( .INP(n1045), .ZN(n1044) );
  INVX0 U1328 ( .INP(n1053), .ZN(n1052) );
  INVX0 U1329 ( .INP(n1061), .ZN(n1060) );
  INVX0 U1330 ( .INP(n1069), .ZN(n1068) );
  INVX0 U1331 ( .INP(n1077), .ZN(n1076) );
  INVX0 U1332 ( .INP(n1085), .ZN(n1084) );
  INVX0 U1333 ( .INP(n1093), .ZN(n1092) );
  INVX0 U1334 ( .INP(n1101), .ZN(n1100) );
  INVX0 U1335 ( .INP(n1109), .ZN(n1108) );
  INVX0 U1336 ( .INP(n1117), .ZN(n1116) );
  INVX0 U1337 ( .INP(n1125), .ZN(n1124) );
  INVX0 U1338 ( .INP(n1133), .ZN(n1132) );
  INVX0 U1339 ( .INP(n1141), .ZN(n1140) );
  INVX0 U1340 ( .INP(n1149), .ZN(n1148) );
  INVX0 U1341 ( .INP(n1157), .ZN(n1156) );
  INVX0 U1342 ( .INP(n1165), .ZN(n1164) );
endmodule


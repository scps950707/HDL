
module pipealu_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447;

  AO21X1 U698 ( .IN1(n1321), .IN2(n1322), .IN3(n1323), .Q(GE_LT_GT_LE) );
  NOR4X0 U699 ( .IN1(n1324), .IN2(n1325), .IN3(n1326), .IN4(n1327), .QN(n1323)
         );
  NAND4X0 U700 ( .IN1(n1328), .IN2(n1329), .IN3(n1419), .IN4(n1330), .QN(n1324) );
  NAND4X0 U703 ( .IN1(n1425), .IN2(n1421), .IN3(n1334), .IN4(n1335), .QN(n1333) );
  OR2X1 U704 ( .IN1(n1443), .IN2(B[8]), .Q(n1335) );
  NAND3X0 U705 ( .IN1(n1338), .IN2(n1339), .IN3(n1332), .QN(n1328) );
  AND2X1 U706 ( .IN1(n1340), .IN2(n1341), .Q(n1332) );
  AO221X1 U707 ( .IN1(n1342), .IN2(n1337), .IN3(n1343), .IN4(n1342), .IN5(
        n1336), .Q(n1341) );
  NAND3X0 U708 ( .IN1(n1344), .IN2(n1345), .IN3(n1422), .QN(n1336) );
  OR2X1 U709 ( .IN1(n1441), .IN2(B[12]), .Q(n1345) );
  NAND3X0 U711 ( .IN1(n1334), .IN2(n1443), .IN3(B[8]), .QN(n1347) );
  AO21X1 U713 ( .IN1(A[10]), .IN2(n1426), .IN3(n1348), .Q(n1337) );
  AOI22X1 U714 ( .IN1(B[11]), .IN2(n1442), .IN3(n1349), .IN4(B[10]), .QN(n1342) );
  AO22X1 U717 ( .IN1(n1350), .IN2(n1351), .IN3(n1351), .IN4(n1346), .Q(n1340)
         );
  AO21X1 U718 ( .IN1(A[14]), .IN2(n1423), .IN3(n1352), .Q(n1346) );
  AOI22X1 U719 ( .IN1(B[15]), .IN2(n1440), .IN3(n1353), .IN4(B[14]), .QN(n1351) );
  NAND3X0 U723 ( .IN1(n1344), .IN2(n1441), .IN3(B[12]), .QN(n1354) );
  AO22X1 U725 ( .IN1(n1355), .IN2(n1356), .IN3(n1356), .IN4(n1357), .Q(n1339)
         );
  AOI22X1 U726 ( .IN1(B[7]), .IN2(n1444), .IN3(n1358), .IN4(B[6]), .QN(n1356)
         );
  NAND3X0 U729 ( .IN1(n1361), .IN2(n1445), .IN3(B[4]), .QN(n1360) );
  NAND3X0 U730 ( .IN1(n1428), .IN2(n1362), .IN3(n1363), .QN(n1338) );
  OA221X1 U731 ( .IN1(n1364), .IN2(n1365), .IN3(B[4]), .IN4(n1445), .IN5(n1361), .Q(n1363) );
  AOI21X1 U733 ( .IN1(n1431), .IN2(A[2]), .IN3(n1366), .QN(n1364) );
  AO221X1 U734 ( .IN1(B[1]), .IN2(n1447), .IN3(n1367), .IN4(B[0]), .IN5(n1365), 
        .Q(n1362) );
  AO22X1 U735 ( .IN1(B[3]), .IN2(n1446), .IN3(n1368), .IN4(B[2]), .Q(n1365) );
  AO21X1 U740 ( .IN1(A[6]), .IN2(n1429), .IN3(n1359), .Q(n1357) );
  NAND4X0 U743 ( .IN1(n1410), .IN2(n1406), .IN3(n1370), .IN4(n1371), .QN(n1327) );
  OR2X1 U744 ( .IN1(n1435), .IN2(B[24]), .Q(n1371) );
  AO221X1 U745 ( .IN1(n1375), .IN2(n1376), .IN3(n1377), .IN4(n1413), .IN5(
        n1374), .Q(n1321) );
  AO221X1 U747 ( .IN1(n1380), .IN2(n1373), .IN3(n1381), .IN4(n1380), .IN5(
        n1372), .Q(n1379) );
  NAND3X0 U748 ( .IN1(n1382), .IN2(n1383), .IN3(n1407), .QN(n1372) );
  OR2X1 U749 ( .IN1(n1433), .IN2(B[28]), .Q(n1383) );
  NAND3X0 U751 ( .IN1(n1370), .IN2(n1435), .IN3(B[24]), .QN(n1385) );
  AO21X1 U753 ( .IN1(A[26]), .IN2(n1411), .IN3(n1386), .Q(n1373) );
  AOI22X1 U754 ( .IN1(B[27]), .IN2(n1434), .IN3(n1387), .IN4(B[26]), .QN(n1380) );
  AO22X1 U757 ( .IN1(n1388), .IN2(n1389), .IN3(n1389), .IN4(n1384), .Q(n1378)
         );
  AO21X1 U758 ( .IN1(A[30]), .IN2(n1408), .IN3(n1390), .Q(n1384) );
  AOI22X1 U759 ( .IN1(B[31]), .IN2(n1432), .IN3(n1391), .IN4(B[30]), .QN(n1389) );
  NAND3X0 U763 ( .IN1(n1382), .IN2(n1433), .IN3(B[28]), .QN(n1392) );
  NAND3X0 U765 ( .IN1(n1415), .IN2(n1393), .IN3(n1394), .QN(n1326) );
  AO221X1 U768 ( .IN1(B[17]), .IN2(n1439), .IN3(n1398), .IN4(B[16]), .IN5(
        n1396), .Q(n1397) );
  AO22X1 U771 ( .IN1(B[19]), .IN2(n1438), .IN3(n1399), .IN4(B[18]), .Q(n1396)
         );
  AO21X1 U773 ( .IN1(A[18]), .IN2(n1418), .IN3(n1400), .Q(n1325) );
  OR2X1 U775 ( .IN1(n1401), .IN2(n1394), .Q(n1376) );
  AOI21X1 U776 ( .IN1(A[22]), .IN2(n1414), .IN3(n1402), .QN(n1394) );
  AO221X1 U777 ( .IN1(B[21]), .IN2(n1437), .IN3(n1403), .IN4(B[20]), .IN5(
        n1401), .Q(n1375) );
  AO22X1 U778 ( .IN1(B[23]), .IN2(n1436), .IN3(n1404), .IN4(B[22]), .Q(n1401)
         );
  INVX0 U655 ( .INP(n1374), .ZN(n1405) );
  INVX0 U656 ( .INP(n1336), .ZN(n1421) );
  INVX0 U657 ( .INP(n1357), .ZN(n1428) );
  NAND2X1 U658 ( .IN1(A[16]), .IN2(n1420), .QN(n1330) );
  INVX0 U659 ( .INP(n1331), .ZN(n1419) );
  NAND2X1 U660 ( .IN1(A[20]), .IN2(n1416), .QN(n1393) );
  INVX0 U661 ( .INP(n1395), .ZN(n1415) );
  INVX0 U662 ( .INP(B[20]), .ZN(n1416) );
  INVX0 U663 ( .INP(n1346), .ZN(n1422) );
  INVX0 U664 ( .INP(n1384), .ZN(n1407) );
  NOR2X0 U665 ( .IN1(n1439), .IN2(B[17]), .QN(n1331) );
  NOR2X0 U666 ( .IN1(n1437), .IN2(B[21]), .QN(n1395) );
  NOR2X0 U667 ( .IN1(n1446), .IN2(B[3]), .QN(n1366) );
  NOR2X0 U668 ( .IN1(n1436), .IN2(B[23]), .QN(n1402) );
  NOR2X0 U669 ( .IN1(n1438), .IN2(B[19]), .QN(n1400) );
  NOR2X0 U670 ( .IN1(n1442), .IN2(B[11]), .QN(n1348) );
  NOR2X0 U671 ( .IN1(n1440), .IN2(B[15]), .QN(n1352) );
  NOR2X0 U672 ( .IN1(n1444), .IN2(B[7]), .QN(n1359) );
  NOR2X0 U673 ( .IN1(n1434), .IN2(B[27]), .QN(n1386) );
  NOR2X0 U674 ( .IN1(n1432), .IN2(B[31]), .QN(n1390) );
  OA21X1 U675 ( .IN1(A[5]), .IN2(n1430), .IN3(n1360), .Q(n1355) );
  INVX0 U676 ( .INP(A[17]), .ZN(n1439) );
  INVX0 U677 ( .INP(A[21]), .ZN(n1437) );
  INVX0 U678 ( .INP(A[3]), .ZN(n1446) );
  INVX0 U679 ( .INP(A[23]), .ZN(n1436) );
  INVX0 U680 ( .INP(A[19]), .ZN(n1438) );
  INVX0 U681 ( .INP(B[18]), .ZN(n1418) );
  INVX0 U682 ( .INP(A[11]), .ZN(n1442) );
  INVX0 U683 ( .INP(A[15]), .ZN(n1440) );
  INVX0 U684 ( .INP(A[7]), .ZN(n1444) );
  INVX0 U685 ( .INP(A[27]), .ZN(n1434) );
  INVX0 U686 ( .INP(A[31]), .ZN(n1432) );
  INVX0 U687 ( .INP(B[9]), .ZN(n1427) );
  INVX0 U688 ( .INP(B[13]), .ZN(n1424) );
  INVX0 U689 ( .INP(B[5]), .ZN(n1430) );
  INVX0 U690 ( .INP(B[25]), .ZN(n1412) );
  INVX0 U691 ( .INP(B[29]), .ZN(n1409) );
  NOR2X0 U692 ( .IN1(A[22]), .IN2(n1402), .QN(n1404) );
  INVX0 U693 ( .INP(B[6]), .ZN(n1429) );
  INVX0 U694 ( .INP(B[14]), .ZN(n1423) );
  INVX0 U695 ( .INP(B[30]), .ZN(n1408) );
  INVX0 U696 ( .INP(B[10]), .ZN(n1426) );
  INVX0 U697 ( .INP(B[26]), .ZN(n1411) );
  NOR2X0 U701 ( .IN1(A[0]), .IN2(n1369), .QN(n1367) );
  NOR2X0 U702 ( .IN1(B[1]), .IN2(n1447), .QN(n1369) );
  INVX0 U710 ( .INP(A[1]), .ZN(n1447) );
  OA21X1 U712 ( .IN1(A[13]), .IN2(n1424), .IN3(n1354), .Q(n1350) );
  NOR2X0 U715 ( .IN1(A[16]), .IN2(n1331), .QN(n1398) );
  NOR2X0 U716 ( .IN1(A[20]), .IN2(n1395), .QN(n1403) );
  NOR2X0 U720 ( .IN1(A[2]), .IN2(n1366), .QN(n1368) );
  INVX0 U721 ( .INP(n1326), .ZN(n1413) );
  NOR2X0 U722 ( .IN1(A[18]), .IN2(n1400), .QN(n1399) );
  INVX0 U724 ( .INP(A[12]), .ZN(n1441) );
  INVX0 U727 ( .INP(A[8]), .ZN(n1443) );
  INVX0 U728 ( .INP(A[28]), .ZN(n1433) );
  INVX0 U732 ( .INP(A[24]), .ZN(n1435) );
  NAND2X1 U736 ( .IN1(A[13]), .IN2(n1424), .QN(n1344) );
  NAND2X1 U737 ( .IN1(A[29]), .IN2(n1409), .QN(n1382) );
  NAND2X1 U738 ( .IN1(A[9]), .IN2(n1427), .QN(n1334) );
  NAND2X1 U739 ( .IN1(A[25]), .IN2(n1412), .QN(n1370) );
  INVX0 U741 ( .INP(B[16]), .ZN(n1420) );
  NAND2X1 U742 ( .IN1(A[5]), .IN2(n1430), .QN(n1361) );
  INVX0 U746 ( .INP(A[4]), .ZN(n1445) );
  NAND2X1 U750 ( .IN1(n1378), .IN2(n1379), .QN(n1374) );
  OA21X1 U752 ( .IN1(A[29]), .IN2(n1409), .IN3(n1392), .Q(n1388) );
  INVX0 U755 ( .INP(B[2]), .ZN(n1431) );
  NAND2X1 U756 ( .IN1(n1332), .IN2(n1333), .QN(n1329) );
  INVX0 U760 ( .INP(n1337), .ZN(n1425) );
  OA21X1 U761 ( .IN1(A[9]), .IN2(n1427), .IN3(n1347), .Q(n1343) );
  OA21X1 U762 ( .IN1(A[25]), .IN2(n1412), .IN3(n1385), .Q(n1381) );
  NAND2X1 U764 ( .IN1(n1405), .IN2(n1327), .QN(n1322) );
  OA21X1 U766 ( .IN1(n1417), .IN2(n1396), .IN3(n1397), .Q(n1377) );
  INVX0 U767 ( .INP(n1325), .ZN(n1417) );
  NOR2X0 U769 ( .IN1(A[10]), .IN2(n1348), .QN(n1349) );
  NOR2X0 U770 ( .IN1(A[26]), .IN2(n1386), .QN(n1387) );
  INVX0 U772 ( .INP(B[22]), .ZN(n1414) );
  NOR2X0 U774 ( .IN1(A[14]), .IN2(n1352), .QN(n1353) );
  NOR2X0 U779 ( .IN1(A[6]), .IN2(n1359), .QN(n1358) );
  NOR2X0 U780 ( .IN1(A[30]), .IN2(n1390), .QN(n1391) );
  INVX0 U781 ( .INP(n1373), .ZN(n1410) );
  INVX0 U782 ( .INP(n1372), .ZN(n1406) );
endmodule


module pipealu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] DIFF;
  input CI;
  output CO;
  wire   n70, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69;
  wire   [33:0] carry;

  FADDX1 U2_31 ( .A(A[31]), .B(n37), .CI(carry[31]), .CO(carry[32]), .S(
        DIFF[31]) );
  FADDX1 U2_30 ( .A(A[30]), .B(n38), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  FADDX1 U2_29 ( .A(A[29]), .B(n39), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  FADDX1 U2_28 ( .A(A[28]), .B(n40), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  FADDX1 U2_27 ( .A(A[27]), .B(n41), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  FADDX1 U2_26 ( .A(A[26]), .B(n42), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  FADDX1 U2_25 ( .A(A[25]), .B(n43), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  FADDX1 U2_24 ( .A(A[24]), .B(n44), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  FADDX1 U2_23 ( .A(A[23]), .B(n45), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1 U2_22 ( .A(A[22]), .B(n46), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n47), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n48), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n49), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n50), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n51), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n52), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n53), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n54), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n55), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n56), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n57), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n58), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n59), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n60), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_7 ( .A(A[7]), .B(n61), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  FADDX1 U2_6 ( .A(A[6]), .B(n62), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FADDX1 U2_5 ( .A(A[5]), .B(n63), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  FADDX1 U2_4 ( .A(A[4]), .B(n64), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  FADDX1 U2_3 ( .A(A[3]), .B(n65), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n66), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n67), .CI(n68), .CO(carry[2]), .S(DIFF[1]) );
  AO21X1 U36 ( .IN1(A[0]), .IN2(n69), .IN3(n70), .Q(DIFF[0]) );
  INVX0 U1 ( .INP(carry[32]), .ZN(DIFF[32]) );
  INVX0 U2 ( .INP(B[16]), .ZN(n52) );
  INVX0 U3 ( .INP(B[20]), .ZN(n48) );
  INVX0 U4 ( .INP(B[6]), .ZN(n62) );
  INVX0 U5 ( .INP(B[10]), .ZN(n58) );
  INVX0 U6 ( .INP(B[14]), .ZN(n54) );
  INVX0 U7 ( .INP(B[18]), .ZN(n50) );
  INVX0 U8 ( .INP(B[26]), .ZN(n42) );
  INVX0 U9 ( .INP(B[30]), .ZN(n38) );
  INVX0 U10 ( .INP(B[5]), .ZN(n63) );
  INVX0 U11 ( .INP(B[9]), .ZN(n59) );
  INVX0 U12 ( .INP(B[13]), .ZN(n55) );
  INVX0 U13 ( .INP(B[25]), .ZN(n43) );
  INVX0 U14 ( .INP(B[29]), .ZN(n39) );
  INVX0 U15 ( .INP(B[22]), .ZN(n46) );
  INVX0 U16 ( .INP(B[2]), .ZN(n66) );
  INVX0 U17 ( .INP(B[1]), .ZN(n67) );
  INVX0 U18 ( .INP(n70), .ZN(n68) );
  INVX0 U19 ( .INP(B[3]), .ZN(n65) );
  INVX0 U20 ( .INP(B[4]), .ZN(n64) );
  INVX0 U21 ( .INP(B[7]), .ZN(n61) );
  INVX0 U22 ( .INP(B[8]), .ZN(n60) );
  INVX0 U23 ( .INP(B[11]), .ZN(n57) );
  INVX0 U24 ( .INP(B[12]), .ZN(n56) );
  INVX0 U25 ( .INP(B[15]), .ZN(n53) );
  INVX0 U26 ( .INP(B[17]), .ZN(n51) );
  INVX0 U27 ( .INP(B[19]), .ZN(n49) );
  INVX0 U28 ( .INP(B[21]), .ZN(n47) );
  INVX0 U29 ( .INP(B[23]), .ZN(n45) );
  INVX0 U30 ( .INP(B[24]), .ZN(n44) );
  INVX0 U31 ( .INP(B[27]), .ZN(n41) );
  INVX0 U32 ( .INP(B[28]), .ZN(n40) );
  NOR2X0 U33 ( .IN1(n69), .IN2(A[0]), .QN(n70) );
  INVX0 U34 ( .INP(B[31]), .ZN(n37) );
  INVX0 U35 ( .INP(B[0]), .ZN(n69) );
endmodule


module pipealu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [32:1] carry;

  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(SUM[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module pipealu ( instr, AluOut, Zero, clk, Carryout, Overflow, rst );
  input [15:0] instr;
  output [31:0] AluOut;
  input clk, rst;
  output Zero, Carryout, Overflow;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, \regfile[15][31] ,
         \regfile[15][30] , \regfile[15][29] , \regfile[15][28] ,
         \regfile[15][27] , \regfile[15][26] , \regfile[15][25] ,
         \regfile[15][24] , \regfile[15][23] , \regfile[15][22] ,
         \regfile[15][21] , \regfile[15][20] , \regfile[15][19] ,
         \regfile[15][18] , \regfile[15][17] , \regfile[15][16] ,
         \regfile[15][15] , \regfile[15][14] , \regfile[15][13] ,
         \regfile[15][12] , \regfile[15][11] , \regfile[15][10] ,
         \regfile[15][9] , \regfile[15][8] , \regfile[15][7] ,
         \regfile[15][6] , \regfile[15][5] , \regfile[15][4] ,
         \regfile[15][3] , \regfile[15][2] , \regfile[15][1] ,
         \regfile[15][0] , \regfile[14][31] , \regfile[14][30] ,
         \regfile[14][29] , \regfile[14][28] , \regfile[14][27] ,
         \regfile[14][26] , \regfile[14][25] , \regfile[14][24] ,
         \regfile[14][23] , \regfile[14][22] , \regfile[14][21] ,
         \regfile[14][20] , \regfile[14][19] , \regfile[14][18] ,
         \regfile[14][17] , \regfile[14][16] , \regfile[14][15] ,
         \regfile[14][14] , \regfile[14][13] , \regfile[14][12] ,
         \regfile[14][11] , \regfile[14][10] , \regfile[14][9] ,
         \regfile[14][8] , \regfile[14][7] , \regfile[14][6] ,
         \regfile[14][5] , \regfile[14][4] , \regfile[14][3] ,
         \regfile[14][2] , \regfile[14][1] , \regfile[14][0] ,
         \regfile[13][31] , \regfile[13][30] , \regfile[13][29] ,
         \regfile[13][28] , \regfile[13][27] , \regfile[13][26] ,
         \regfile[13][25] , \regfile[13][24] , \regfile[13][23] ,
         \regfile[13][22] , \regfile[13][21] , \regfile[13][20] ,
         \regfile[13][19] , \regfile[13][18] , \regfile[13][17] ,
         \regfile[13][16] , \regfile[13][15] , \regfile[13][14] ,
         \regfile[13][13] , \regfile[13][12] , \regfile[13][11] ,
         \regfile[13][10] , \regfile[13][9] , \regfile[13][8] ,
         \regfile[13][7] , \regfile[13][6] , \regfile[13][5] ,
         \regfile[13][4] , \regfile[13][3] , \regfile[13][2] ,
         \regfile[13][1] , \regfile[13][0] , \regfile[12][31] ,
         \regfile[12][30] , \regfile[12][29] , \regfile[12][28] ,
         \regfile[12][27] , \regfile[12][26] , \regfile[12][25] ,
         \regfile[12][24] , \regfile[12][23] , \regfile[12][22] ,
         \regfile[12][21] , \regfile[12][20] , \regfile[12][19] ,
         \regfile[12][18] , \regfile[12][17] , \regfile[12][16] ,
         \regfile[12][15] , \regfile[12][14] , \regfile[12][13] ,
         \regfile[12][12] , \regfile[12][11] , \regfile[12][10] ,
         \regfile[12][9] , \regfile[12][8] , \regfile[12][7] ,
         \regfile[12][6] , \regfile[12][5] , \regfile[12][4] ,
         \regfile[12][3] , \regfile[12][2] , \regfile[12][1] ,
         \regfile[12][0] , \regfile[11][31] , \regfile[11][30] ,
         \regfile[11][29] , \regfile[11][28] , \regfile[11][27] ,
         \regfile[11][26] , \regfile[11][25] , \regfile[11][24] ,
         \regfile[11][23] , \regfile[11][22] , \regfile[11][21] ,
         \regfile[11][20] , \regfile[11][19] , \regfile[11][18] ,
         \regfile[11][17] , \regfile[11][16] , \regfile[11][15] ,
         \regfile[11][14] , \regfile[11][13] , \regfile[11][12] ,
         \regfile[11][11] , \regfile[11][10] , \regfile[11][9] ,
         \regfile[11][8] , \regfile[11][7] , \regfile[11][6] ,
         \regfile[11][5] , \regfile[11][4] , \regfile[11][3] ,
         \regfile[11][2] , \regfile[11][1] , \regfile[11][0] ,
         \regfile[10][31] , \regfile[10][30] , \regfile[10][29] ,
         \regfile[10][28] , \regfile[10][27] , \regfile[10][26] ,
         \regfile[10][25] , \regfile[10][24] , \regfile[10][23] ,
         \regfile[10][22] , \regfile[10][21] , \regfile[10][20] ,
         \regfile[10][19] , \regfile[10][18] , \regfile[10][17] ,
         \regfile[10][16] , \regfile[10][15] , \regfile[10][14] ,
         \regfile[10][13] , \regfile[10][12] , \regfile[10][11] ,
         \regfile[10][10] , \regfile[10][9] , \regfile[10][8] ,
         \regfile[10][7] , \regfile[10][6] , \regfile[10][5] ,
         \regfile[10][4] , \regfile[10][3] , \regfile[10][2] ,
         \regfile[10][1] , \regfile[10][0] , \regfile[9][31] ,
         \regfile[9][30] , \regfile[9][29] , \regfile[9][28] ,
         \regfile[9][27] , \regfile[9][26] , \regfile[9][25] ,
         \regfile[9][24] , \regfile[9][23] , \regfile[9][22] ,
         \regfile[9][21] , \regfile[9][20] , \regfile[9][19] ,
         \regfile[9][18] , \regfile[9][17] , \regfile[9][16] ,
         \regfile[9][15] , \regfile[9][14] , \regfile[9][13] ,
         \regfile[9][12] , \regfile[9][11] , \regfile[9][10] , \regfile[9][9] ,
         \regfile[9][8] , \regfile[9][7] , \regfile[9][6] , \regfile[9][5] ,
         \regfile[9][4] , \regfile[9][3] , \regfile[9][2] , \regfile[9][1] ,
         \regfile[9][0] , \regfile[8][31] , \regfile[8][30] , \regfile[8][29] ,
         \regfile[8][28] , \regfile[8][27] , \regfile[8][26] ,
         \regfile[8][25] , \regfile[8][24] , \regfile[8][23] ,
         \regfile[8][22] , \regfile[8][21] , \regfile[8][20] ,
         \regfile[8][19] , \regfile[8][18] , \regfile[8][17] ,
         \regfile[8][16] , \regfile[8][15] , \regfile[8][14] ,
         \regfile[8][13] , \regfile[8][12] , \regfile[8][11] ,
         \regfile[8][10] , \regfile[8][9] , \regfile[8][8] , \regfile[8][7] ,
         \regfile[8][6] , \regfile[8][5] , \regfile[8][4] , \regfile[8][3] ,
         \regfile[8][2] , \regfile[8][1] , \regfile[8][0] , \regfile[7][31] ,
         \regfile[7][30] , \regfile[7][29] , \regfile[7][28] ,
         \regfile[7][27] , \regfile[7][26] , \regfile[7][25] ,
         \regfile[7][24] , \regfile[7][23] , \regfile[7][22] ,
         \regfile[7][21] , \regfile[7][20] , \regfile[7][19] ,
         \regfile[7][18] , \regfile[7][17] , \regfile[7][16] ,
         \regfile[7][15] , \regfile[7][14] , \regfile[7][13] ,
         \regfile[7][12] , \regfile[7][11] , \regfile[7][10] , \regfile[7][9] ,
         \regfile[7][8] , \regfile[7][7] , \regfile[7][6] , \regfile[7][5] ,
         \regfile[7][4] , \regfile[7][3] , \regfile[7][2] , \regfile[7][1] ,
         \regfile[7][0] , \regfile[6][31] , \regfile[6][30] , \regfile[6][29] ,
         \regfile[6][28] , \regfile[6][27] , \regfile[6][26] ,
         \regfile[6][25] , \regfile[6][24] , \regfile[6][23] ,
         \regfile[6][22] , \regfile[6][21] , \regfile[6][20] ,
         \regfile[6][19] , \regfile[6][18] , \regfile[6][17] ,
         \regfile[6][16] , \regfile[6][15] , \regfile[6][14] ,
         \regfile[6][13] , \regfile[6][12] , \regfile[6][11] ,
         \regfile[6][10] , \regfile[6][9] , \regfile[6][8] , \regfile[6][7] ,
         \regfile[6][6] , \regfile[6][5] , \regfile[6][4] , \regfile[6][3] ,
         \regfile[6][2] , \regfile[6][1] , \regfile[6][0] , \regfile[5][31] ,
         \regfile[5][30] , \regfile[5][29] , \regfile[5][28] ,
         \regfile[5][27] , \regfile[5][26] , \regfile[5][25] ,
         \regfile[5][24] , \regfile[5][23] , \regfile[5][22] ,
         \regfile[5][21] , \regfile[5][20] , \regfile[5][19] ,
         \regfile[5][18] , \regfile[5][17] , \regfile[5][16] ,
         \regfile[5][15] , \regfile[5][14] , \regfile[5][13] ,
         \regfile[5][12] , \regfile[5][11] , \regfile[5][10] , \regfile[5][9] ,
         \regfile[5][8] , \regfile[5][7] , \regfile[5][6] , \regfile[5][5] ,
         \regfile[5][4] , \regfile[5][3] , \regfile[5][2] , \regfile[5][1] ,
         \regfile[5][0] , \regfile[4][31] , \regfile[4][30] , \regfile[4][29] ,
         \regfile[4][28] , \regfile[4][27] , \regfile[4][26] ,
         \regfile[4][25] , \regfile[4][24] , \regfile[4][23] ,
         \regfile[4][22] , \regfile[4][21] , \regfile[4][20] ,
         \regfile[4][19] , \regfile[4][18] , \regfile[4][17] ,
         \regfile[4][16] , \regfile[4][15] , \regfile[4][14] ,
         \regfile[4][13] , \regfile[4][12] , \regfile[4][11] ,
         \regfile[4][10] , \regfile[4][9] , \regfile[4][8] , \regfile[4][7] ,
         \regfile[4][6] , \regfile[4][5] , \regfile[4][4] , \regfile[4][3] ,
         \regfile[4][2] , \regfile[4][1] , \regfile[4][0] , \regfile[3][31] ,
         \regfile[3][30] , \regfile[3][29] , \regfile[3][28] ,
         \regfile[3][27] , \regfile[3][26] , \regfile[3][25] ,
         \regfile[3][24] , \regfile[3][23] , \regfile[3][22] ,
         \regfile[3][21] , \regfile[3][20] , \regfile[3][19] ,
         \regfile[3][18] , \regfile[3][17] , \regfile[3][16] ,
         \regfile[3][15] , \regfile[3][14] , \regfile[3][13] ,
         \regfile[3][12] , \regfile[3][11] , \regfile[3][10] , \regfile[3][9] ,
         \regfile[3][8] , \regfile[3][7] , \regfile[3][6] , \regfile[3][5] ,
         \regfile[3][4] , \regfile[3][3] , \regfile[3][2] , \regfile[3][1] ,
         \regfile[3][0] , \regfile[2][31] , \regfile[2][30] , \regfile[2][29] ,
         \regfile[2][28] , \regfile[2][27] , \regfile[2][26] ,
         \regfile[2][25] , \regfile[2][24] , \regfile[2][23] ,
         \regfile[2][22] , \regfile[2][21] , \regfile[2][20] ,
         \regfile[2][19] , \regfile[2][18] , \regfile[2][17] ,
         \regfile[2][16] , \regfile[2][15] , \regfile[2][14] ,
         \regfile[2][13] , \regfile[2][12] , \regfile[2][11] ,
         \regfile[2][10] , \regfile[2][9] , \regfile[2][8] , \regfile[2][7] ,
         \regfile[2][6] , \regfile[2][5] , \regfile[2][4] , \regfile[2][3] ,
         \regfile[2][2] , \regfile[2][1] , \regfile[2][0] , \regfile[1][31] ,
         \regfile[1][30] , \regfile[1][29] , \regfile[1][28] ,
         \regfile[1][27] , \regfile[1][26] , \regfile[1][25] ,
         \regfile[1][24] , \regfile[1][23] , \regfile[1][22] ,
         \regfile[1][21] , \regfile[1][20] , \regfile[1][19] ,
         \regfile[1][18] , \regfile[1][17] , \regfile[1][16] ,
         \regfile[1][15] , \regfile[1][14] , \regfile[1][13] ,
         \regfile[1][12] , \regfile[1][11] , \regfile[1][10] , \regfile[1][9] ,
         \regfile[1][8] , \regfile[1][7] , \regfile[1][6] , \regfile[1][5] ,
         \regfile[1][4] , \regfile[1][3] , \regfile[1][2] , \regfile[1][1] ,
         \regfile[1][0] , \regfile[0][31] , \regfile[0][30] , \regfile[0][29] ,
         \regfile[0][28] , \regfile[0][27] , \regfile[0][26] ,
         \regfile[0][25] , \regfile[0][24] , \regfile[0][23] ,
         \regfile[0][22] , \regfile[0][21] , \regfile[0][20] ,
         \regfile[0][19] , \regfile[0][18] , \regfile[0][17] ,
         \regfile[0][16] , \regfile[0][15] , \regfile[0][14] ,
         \regfile[0][13] , \regfile[0][12] , \regfile[0][11] ,
         \regfile[0][10] , \regfile[0][9] , \regfile[0][8] , \regfile[0][7] ,
         \regfile[0][6] , \regfile[0][5] , \regfile[0][4] , \regfile[0][3] ,
         \regfile[0][2] , \regfile[0][1] , \regfile[0][0] , N191, N192, N193,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N259, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n966, n967, n968,
         n969, n970, n971, n972, n973, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853;
  wire   [31:0] IFID_A;
  wire   [31:0] IFID_B;
  wire   [3:0] IFID_dest;
  assign N17 = instr[8];
  assign N18 = instr[9];
  assign N19 = instr[10];
  assign N20 = instr[11];
  assign N21 = instr[4];
  assign N22 = instr[5];
  assign N23 = instr[6];
  assign N24 = instr[7];

  DFFX1 Carryout_reg ( .D(N324), .CLK(clk), .Q(Carryout) );
  DFFX1 \EX_dest_reg[3]  ( .D(IFID_dest[3]), .CLK(clk), .Q(n967) );
  DFFX1 \EX_dest_reg[2]  ( .D(IFID_dest[2]), .CLK(clk), .Q(n970) );
  DFFX1 \EX_dest_reg[1]  ( .D(IFID_dest[1]), .CLK(clk), .Q(n969), .QN(n3224)
         );
  DFFX1 \EX_dest_reg[0]  ( .D(IFID_dest[0]), .CLK(clk), .Q(n968), .QN(n3225)
         );
  DFFX1 Overflow_reg ( .D(N325), .CLK(clk), .Q(Overflow) );
  DFFX1 \AluOut_reg[31]  ( .D(N323), .CLK(clk), .Q(AluOut[31]), .QN(n312) );
  DFFX1 \AluOut_reg[30]  ( .D(N322), .CLK(clk), .Q(AluOut[30]), .QN(n307) );
  DFFX1 \AluOut_reg[29]  ( .D(N321), .CLK(clk), .Q(AluOut[29]), .QN(n306) );
  DFFX1 \AluOut_reg[28]  ( .D(N320), .CLK(clk), .Q(AluOut[28]), .QN(n305) );
  DFFX1 \AluOut_reg[27]  ( .D(N319), .CLK(clk), .Q(AluOut[27]), .QN(n304) );
  DFFX1 \AluOut_reg[26]  ( .D(N318), .CLK(clk), .Q(AluOut[26]), .QN(n303) );
  DFFX1 \AluOut_reg[25]  ( .D(N317), .CLK(clk), .Q(AluOut[25]), .QN(n302) );
  DFFX1 \AluOut_reg[24]  ( .D(N316), .CLK(clk), .Q(AluOut[24]), .QN(n301) );
  DFFX1 \AluOut_reg[23]  ( .D(N315), .CLK(clk), .Q(AluOut[23]), .QN(n300) );
  DFFX1 \AluOut_reg[22]  ( .D(N314), .CLK(clk), .Q(AluOut[22]), .QN(n299) );
  DFFX1 \AluOut_reg[21]  ( .D(N313), .CLK(clk), .Q(AluOut[21]), .QN(n298) );
  DFFX1 \AluOut_reg[20]  ( .D(N312), .CLK(clk), .Q(AluOut[20]), .QN(n297) );
  DFFX1 \AluOut_reg[19]  ( .D(N311), .CLK(clk), .Q(AluOut[19]), .QN(n296) );
  DFFX1 \AluOut_reg[18]  ( .D(N310), .CLK(clk), .Q(AluOut[18]), .QN(n295) );
  DFFX1 \AluOut_reg[17]  ( .D(N309), .CLK(clk), .Q(AluOut[17]), .QN(n294) );
  DFFX1 \AluOut_reg[16]  ( .D(N308), .CLK(clk), .Q(AluOut[16]), .QN(n293) );
  DFFX1 \AluOut_reg[15]  ( .D(N307), .CLK(clk), .Q(AluOut[15]), .QN(n292) );
  DFFX1 \AluOut_reg[14]  ( .D(N306), .CLK(clk), .Q(AluOut[14]), .QN(n291) );
  DFFX1 \AluOut_reg[13]  ( .D(N305), .CLK(clk), .Q(AluOut[13]), .QN(n290) );
  DFFX1 \AluOut_reg[12]  ( .D(N304), .CLK(clk), .Q(AluOut[12]), .QN(n289) );
  DFFX1 \AluOut_reg[11]  ( .D(N303), .CLK(clk), .Q(AluOut[11]), .QN(n288) );
  DFFX1 \AluOut_reg[10]  ( .D(N302), .CLK(clk), .Q(AluOut[10]), .QN(n287) );
  DFFX1 \AluOut_reg[9]  ( .D(N301), .CLK(clk), .Q(AluOut[9]), .QN(n286) );
  DFFX1 \AluOut_reg[8]  ( .D(N300), .CLK(clk), .Q(AluOut[8]), .QN(n285) );
  DFFX1 \AluOut_reg[7]  ( .D(N299), .CLK(clk), .Q(AluOut[7]), .QN(n284) );
  DFFX1 \AluOut_reg[6]  ( .D(N298), .CLK(clk), .Q(AluOut[6]), .QN(n283) );
  DFFX1 \AluOut_reg[5]  ( .D(N297), .CLK(clk), .Q(AluOut[5]), .QN(n282) );
  DFFX1 \AluOut_reg[4]  ( .D(N296), .CLK(clk), .Q(AluOut[4]), .QN(n281) );
  DFFX1 \AluOut_reg[3]  ( .D(N295), .CLK(clk), .Q(AluOut[3]), .QN(n280) );
  DFFX1 \AluOut_reg[2]  ( .D(N294), .CLK(clk), .Q(AluOut[2]), .QN(n279) );
  DFFX1 \AluOut_reg[1]  ( .D(N293), .CLK(clk), .Q(AluOut[1]), .QN(n278) );
  DFFX1 \AluOut_reg[0]  ( .D(N292), .CLK(clk), .Q(AluOut[0]), .QN(n277) );
  DFFX1 \IFID_B_reg[31]  ( .D(n964), .CLK(clk), .Q(IFID_B[31]), .QN(n380) );
  DFFX1 \IFID_B_reg[30]  ( .D(n963), .CLK(clk), .Q(IFID_B[30]), .QN(n379) );
  DFFX1 \IFID_B_reg[29]  ( .D(n962), .CLK(clk), .Q(IFID_B[29]), .QN(n378) );
  DFFX1 \IFID_B_reg[28]  ( .D(n961), .CLK(clk), .Q(IFID_B[28]), .QN(n377) );
  DFFX1 \IFID_B_reg[27]  ( .D(n960), .CLK(clk), .Q(IFID_B[27]), .QN(n376) );
  DFFX1 \IFID_B_reg[26]  ( .D(n959), .CLK(clk), .Q(IFID_B[26]), .QN(n375) );
  DFFX1 \IFID_B_reg[25]  ( .D(n958), .CLK(clk), .Q(IFID_B[25]), .QN(n374) );
  DFFX1 \IFID_B_reg[24]  ( .D(n957), .CLK(clk), .Q(IFID_B[24]), .QN(n373) );
  DFFX1 \IFID_B_reg[23]  ( .D(n956), .CLK(clk), .Q(IFID_B[23]), .QN(n372) );
  DFFX1 \IFID_B_reg[22]  ( .D(n955), .CLK(clk), .Q(IFID_B[22]), .QN(n371) );
  DFFX1 \IFID_B_reg[21]  ( .D(n954), .CLK(clk), .Q(IFID_B[21]), .QN(n370) );
  DFFX1 \IFID_B_reg[20]  ( .D(n953), .CLK(clk), .Q(IFID_B[20]), .QN(n369) );
  DFFX1 \IFID_B_reg[19]  ( .D(n952), .CLK(clk), .Q(IFID_B[19]), .QN(n368) );
  DFFX1 \IFID_B_reg[18]  ( .D(n951), .CLK(clk), .Q(IFID_B[18]), .QN(n367) );
  DFFX1 \IFID_B_reg[17]  ( .D(n950), .CLK(clk), .Q(IFID_B[17]), .QN(n366) );
  DFFX1 \IFID_B_reg[16]  ( .D(n949), .CLK(clk), .Q(IFID_B[16]), .QN(n365) );
  DFFX1 \IFID_B_reg[15]  ( .D(n948), .CLK(clk), .Q(IFID_B[15]), .QN(n364) );
  DFFX1 \IFID_B_reg[14]  ( .D(n947), .CLK(clk), .Q(IFID_B[14]), .QN(n363) );
  DFFX1 \IFID_B_reg[13]  ( .D(n946), .CLK(clk), .Q(IFID_B[13]), .QN(n362) );
  DFFX1 \IFID_B_reg[12]  ( .D(n945), .CLK(clk), .Q(IFID_B[12]), .QN(n361) );
  DFFX1 \IFID_B_reg[11]  ( .D(n944), .CLK(clk), .Q(IFID_B[11]), .QN(n360) );
  DFFX1 \IFID_B_reg[10]  ( .D(n943), .CLK(clk), .Q(IFID_B[10]), .QN(n359) );
  DFFX1 \IFID_B_reg[9]  ( .D(n942), .CLK(clk), .Q(IFID_B[9]), .QN(n358) );
  DFFX1 \IFID_B_reg[8]  ( .D(n941), .CLK(clk), .Q(IFID_B[8]), .QN(n357) );
  DFFX1 \IFID_B_reg[7]  ( .D(n940), .CLK(clk), .Q(IFID_B[7]), .QN(n356) );
  DFFX1 \IFID_B_reg[6]  ( .D(n939), .CLK(clk), .Q(IFID_B[6]), .QN(n355) );
  DFFX1 \IFID_B_reg[5]  ( .D(n938), .CLK(clk), .Q(IFID_B[5]), .QN(n354) );
  DFFX1 \IFID_B_reg[4]  ( .D(n937), .CLK(clk), .Q(IFID_B[4]), .QN(n353) );
  DFFX1 \IFID_B_reg[3]  ( .D(n936), .CLK(clk), .Q(IFID_B[3]), .QN(n352) );
  DFFX1 \IFID_B_reg[2]  ( .D(n935), .CLK(clk), .Q(IFID_B[2]), .QN(n351) );
  DFFX1 \IFID_B_reg[1]  ( .D(n934), .CLK(clk), .Q(IFID_B[1]), .QN(n350) );
  DFFX1 \IFID_B_reg[0]  ( .D(n933), .CLK(clk), .Q(IFID_B[0]), .QN(n349) );
  DFFX1 \IFID_ALU_ctl_reg[3]  ( .D(n932), .CLK(clk), .Q(n972) );
  DFFX1 \IFID_ALU_ctl_reg[2]  ( .D(n931), .CLK(clk), .Q(n966), .QN(n3223) );
  DFFX1 \IFID_ALU_ctl_reg[1]  ( .D(n930), .CLK(clk), .Q(n973), .QN(n2966) );
  DFFX1 \IFID_ALU_ctl_reg[0]  ( .D(n929), .CLK(clk), .Q(n971), .QN(n3482) );
  DFFX1 \IFID_A_reg[31]  ( .D(n928), .CLK(clk), .Q(IFID_A[31]), .QN(n344) );
  DFFX1 \IFID_A_reg[30]  ( .D(n927), .CLK(clk), .Q(IFID_A[30]), .QN(n343) );
  DFFX1 \IFID_A_reg[29]  ( .D(n926), .CLK(clk), .Q(IFID_A[29]), .QN(n342) );
  DFFX1 \IFID_A_reg[28]  ( .D(n925), .CLK(clk), .Q(IFID_A[28]), .QN(n341) );
  DFFX1 \IFID_A_reg[27]  ( .D(n924), .CLK(clk), .Q(IFID_A[27]), .QN(n340) );
  DFFX1 \IFID_A_reg[26]  ( .D(n923), .CLK(clk), .Q(IFID_A[26]), .QN(n339) );
  DFFX1 \IFID_A_reg[25]  ( .D(n922), .CLK(clk), .Q(IFID_A[25]), .QN(n338) );
  DFFX1 \IFID_A_reg[24]  ( .D(n921), .CLK(clk), .Q(IFID_A[24]), .QN(n337) );
  DFFX1 \IFID_A_reg[23]  ( .D(n920), .CLK(clk), .Q(IFID_A[23]), .QN(n336) );
  DFFX1 \IFID_A_reg[22]  ( .D(n919), .CLK(clk), .Q(IFID_A[22]), .QN(n335) );
  DFFX1 \IFID_A_reg[21]  ( .D(n918), .CLK(clk), .Q(IFID_A[21]), .QN(n334) );
  DFFX1 \IFID_A_reg[20]  ( .D(n917), .CLK(clk), .Q(IFID_A[20]), .QN(n333) );
  DFFX1 \IFID_A_reg[19]  ( .D(n916), .CLK(clk), .Q(IFID_A[19]), .QN(n332) );
  DFFX1 \IFID_A_reg[18]  ( .D(n915), .CLK(clk), .Q(IFID_A[18]), .QN(n331) );
  DFFX1 \IFID_A_reg[17]  ( .D(n914), .CLK(clk), .Q(IFID_A[17]), .QN(n330) );
  DFFX1 \IFID_A_reg[16]  ( .D(n913), .CLK(clk), .Q(IFID_A[16]), .QN(n329) );
  DFFX1 \IFID_A_reg[15]  ( .D(n912), .CLK(clk), .Q(IFID_A[15]), .QN(n328) );
  DFFX1 \IFID_A_reg[14]  ( .D(n911), .CLK(clk), .Q(IFID_A[14]), .QN(n327) );
  DFFX1 \IFID_A_reg[13]  ( .D(n910), .CLK(clk), .Q(IFID_A[13]), .QN(n326) );
  DFFX1 \IFID_A_reg[12]  ( .D(n909), .CLK(clk), .Q(IFID_A[12]), .QN(n325) );
  DFFX1 \IFID_A_reg[11]  ( .D(n908), .CLK(clk), .Q(IFID_A[11]), .QN(n324) );
  DFFX1 \IFID_A_reg[10]  ( .D(n907), .CLK(clk), .Q(IFID_A[10]), .QN(n323) );
  DFFX1 \IFID_A_reg[9]  ( .D(n906), .CLK(clk), .Q(IFID_A[9]), .QN(n322) );
  DFFX1 \IFID_A_reg[8]  ( .D(n905), .CLK(clk), .Q(IFID_A[8]), .QN(n321) );
  DFFX1 \IFID_A_reg[7]  ( .D(n904), .CLK(clk), .Q(IFID_A[7]), .QN(n320) );
  DFFX1 \IFID_A_reg[6]  ( .D(n903), .CLK(clk), .Q(IFID_A[6]), .QN(n319) );
  DFFX1 \IFID_A_reg[5]  ( .D(n902), .CLK(clk), .Q(IFID_A[5]), .QN(n318) );
  DFFX1 \IFID_A_reg[4]  ( .D(n901), .CLK(clk), .Q(IFID_A[4]), .QN(n317) );
  DFFX1 \IFID_A_reg[3]  ( .D(n900), .CLK(clk), .Q(IFID_A[3]), .QN(n316) );
  DFFX1 \IFID_A_reg[2]  ( .D(n899), .CLK(clk), .Q(IFID_A[2]), .QN(n315) );
  DFFX1 \IFID_A_reg[1]  ( .D(n898), .CLK(clk), .Q(IFID_A[1]), .QN(n314) );
  DFFX1 \IFID_A_reg[0]  ( .D(n897), .CLK(clk), .Q(IFID_A[0]), .QN(n313) );
  DFFX1 \IFID_dest_reg[3]  ( .D(n896), .CLK(clk), .Q(IFID_dest[3]) );
  DFFX1 \IFID_dest_reg[2]  ( .D(n895), .CLK(clk), .Q(IFID_dest[2]) );
  DFFX1 \IFID_dest_reg[1]  ( .D(n894), .CLK(clk), .Q(IFID_dest[1]) );
  DFFX1 \IFID_dest_reg[0]  ( .D(n893), .CLK(clk), .Q(IFID_dest[0]) );
  DFFARX1 \regfile_reg[0][31]  ( .D(n892), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[0][31] ), .QN(n3086) );
  DFFARX1 \regfile_reg[1][31]  ( .D(n891), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[1][31] ), .QN(n3345) );
  DFFARX1 \regfile_reg[2][31]  ( .D(n890), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[2][31] ), .QN(n3465) );
  DFFARX1 \regfile_reg[3][31]  ( .D(n889), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[3][31] ), .QN(n3217) );
  DFFARX1 \regfile_reg[4][31]  ( .D(n888), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[4][31] ), .QN(n3085) );
  DFFARX1 \regfile_reg[5][31]  ( .D(n887), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[5][31] ), .QN(n3344) );
  DFFARX1 \regfile_reg[6][31]  ( .D(n886), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[6][31] ), .QN(n3464) );
  DFFARX1 \regfile_reg[7][31]  ( .D(n885), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[7][31] ), .QN(n3216) );
  DFFARX1 \regfile_reg[8][31]  ( .D(n884), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][31] ), .QN(n3084) );
  DFFARX1 \regfile_reg[9][31]  ( .D(n883), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[9][31] ), .QN(n3343) );
  DFFARX1 \regfile_reg[10][31]  ( .D(n882), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[10][31] ), .QN(n3463) );
  DFFARX1 \regfile_reg[11][31]  ( .D(n881), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[11][31] ), .QN(n3215) );
  DFFARX1 \regfile_reg[12][31]  ( .D(n880), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[12][31] ), .QN(n3083) );
  DFFARX1 \regfile_reg[13][31]  ( .D(n879), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][31] ), .QN(n3342) );
  DFFARX1 \regfile_reg[14][31]  ( .D(n878), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[14][31] ), .QN(n3462) );
  DFFARX1 \regfile_reg[15][31]  ( .D(n877), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[15][31] ), .QN(n3214) );
  DFFARX1 \regfile_reg[0][30]  ( .D(n876), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[0][30] ), .QN(n3082) );
  DFFARX1 \regfile_reg[1][30]  ( .D(n875), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[1][30] ), .QN(n3341) );
  DFFARX1 \regfile_reg[2][30]  ( .D(n874), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[2][30] ), .QN(n3461) );
  DFFARX1 \regfile_reg[3][30]  ( .D(n873), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[3][30] ), .QN(n3213) );
  DFFARX1 \regfile_reg[4][30]  ( .D(n872), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][30] ), .QN(n3081) );
  DFFARX1 \regfile_reg[5][30]  ( .D(n871), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[5][30] ), .QN(n3340) );
  DFFARX1 \regfile_reg[6][30]  ( .D(n870), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[6][30] ), .QN(n3460) );
  DFFARX1 \regfile_reg[7][30]  ( .D(n869), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[7][30] ), .QN(n3212) );
  DFFARX1 \regfile_reg[8][30]  ( .D(n868), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[8][30] ), .QN(n3080) );
  DFFARX1 \regfile_reg[9][30]  ( .D(n867), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[9][30] ), .QN(n3339) );
  DFFARX1 \regfile_reg[10][30]  ( .D(n866), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[10][30] ), .QN(n3459) );
  DFFARX1 \regfile_reg[11][30]  ( .D(n865), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[11][30] ), .QN(n3211) );
  DFFARX1 \regfile_reg[12][30]  ( .D(n864), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[12][30] ), .QN(n3079) );
  DFFARX1 \regfile_reg[13][30]  ( .D(n863), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[13][30] ), .QN(n3338) );
  DFFARX1 \regfile_reg[14][30]  ( .D(n862), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[14][30] ), .QN(n3458) );
  DFFARX1 \regfile_reg[15][30]  ( .D(n861), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[15][30] ), .QN(n3210) );
  DFFARX1 \regfile_reg[0][29]  ( .D(n860), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[0][29] ), .QN(n3078) );
  DFFARX1 \regfile_reg[1][29]  ( .D(n859), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[1][29] ), .QN(n3337) );
  DFFARX1 \regfile_reg[2][29]  ( .D(n858), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[2][29] ), .QN(n3457) );
  DFFARX1 \regfile_reg[3][29]  ( .D(n857), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[3][29] ), .QN(n3209) );
  DFFARX1 \regfile_reg[4][29]  ( .D(n856), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][29] ), .QN(n3077) );
  DFFARX1 \regfile_reg[5][29]  ( .D(n855), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][29] ), .QN(n3336) );
  DFFARX1 \regfile_reg[6][29]  ( .D(n854), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[6][29] ), .QN(n3456) );
  DFFARX1 \regfile_reg[7][29]  ( .D(n853), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][29] ), .QN(n3208) );
  DFFARX1 \regfile_reg[8][29]  ( .D(n852), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][29] ), .QN(n3076) );
  DFFARX1 \regfile_reg[9][29]  ( .D(n851), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[9][29] ), .QN(n3335) );
  DFFARX1 \regfile_reg[10][29]  ( .D(n850), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[10][29] ), .QN(n3455) );
  DFFARX1 \regfile_reg[11][29]  ( .D(n849), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[11][29] ), .QN(n3207) );
  DFFARX1 \regfile_reg[12][29]  ( .D(n848), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[12][29] ), .QN(n3075) );
  DFFARX1 \regfile_reg[13][29]  ( .D(n847), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[13][29] ), .QN(n3334) );
  DFFARX1 \regfile_reg[14][29]  ( .D(n846), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[14][29] ), .QN(n3454) );
  DFFARX1 \regfile_reg[15][29]  ( .D(n845), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[15][29] ), .QN(n3206) );
  DFFARX1 \regfile_reg[0][28]  ( .D(n844), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][28] ), .QN(n3074) );
  DFFARX1 \regfile_reg[1][28]  ( .D(n843), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][28] ), .QN(n3333) );
  DFFARX1 \regfile_reg[2][28]  ( .D(n842), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[2][28] ), .QN(n3453) );
  DFFARX1 \regfile_reg[3][28]  ( .D(n841), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[3][28] ), .QN(n3205) );
  DFFARX1 \regfile_reg[4][28]  ( .D(n840), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[4][28] ), .QN(n3073) );
  DFFARX1 \regfile_reg[5][28]  ( .D(n839), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[5][28] ), .QN(n3332) );
  DFFARX1 \regfile_reg[6][28]  ( .D(n838), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[6][28] ), .QN(n3452) );
  DFFARX1 \regfile_reg[7][28]  ( .D(n837), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[7][28] ), .QN(n3204) );
  DFFARX1 \regfile_reg[8][28]  ( .D(n836), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[8][28] ), .QN(n3072) );
  DFFARX1 \regfile_reg[9][28]  ( .D(n835), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[9][28] ), .QN(n3331) );
  DFFARX1 \regfile_reg[10][28]  ( .D(n834), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[10][28] ), .QN(n3451) );
  DFFARX1 \regfile_reg[11][28]  ( .D(n833), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[11][28] ), .QN(n3203) );
  DFFARX1 \regfile_reg[12][28]  ( .D(n832), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[12][28] ), .QN(n3071) );
  DFFARX1 \regfile_reg[13][28]  ( .D(n831), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[13][28] ), .QN(n3330) );
  DFFARX1 \regfile_reg[14][28]  ( .D(n830), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[14][28] ), .QN(n3450) );
  DFFARX1 \regfile_reg[15][28]  ( .D(n829), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[15][28] ), .QN(n3202) );
  DFFARX1 \regfile_reg[0][27]  ( .D(n828), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[0][27] ), .QN(n3070) );
  DFFARX1 \regfile_reg[1][27]  ( .D(n827), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[1][27] ), .QN(n3329) );
  DFFARX1 \regfile_reg[2][27]  ( .D(n826), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[2][27] ), .QN(n3449) );
  DFFARX1 \regfile_reg[3][27]  ( .D(n825), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[3][27] ), .QN(n3201) );
  DFFARX1 \regfile_reg[4][27]  ( .D(n824), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][27] ), .QN(n3069) );
  DFFARX1 \regfile_reg[5][27]  ( .D(n823), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][27] ), .QN(n3328) );
  DFFARX1 \regfile_reg[6][27]  ( .D(n822), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[6][27] ), .QN(n3448) );
  DFFARX1 \regfile_reg[7][27]  ( .D(n821), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][27] ), .QN(n3200) );
  DFFARX1 \regfile_reg[8][27]  ( .D(n820), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][27] ), .QN(n3068) );
  DFFARX1 \regfile_reg[9][27]  ( .D(n819), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[9][27] ), .QN(n3327) );
  DFFARX1 \regfile_reg[10][27]  ( .D(n818), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[10][27] ), .QN(n3447) );
  DFFARX1 \regfile_reg[11][27]  ( .D(n817), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[11][27] ), .QN(n3199) );
  DFFARX1 \regfile_reg[12][27]  ( .D(n816), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[12][27] ), .QN(n3067) );
  DFFARX1 \regfile_reg[13][27]  ( .D(n815), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[13][27] ), .QN(n3326) );
  DFFARX1 \regfile_reg[14][27]  ( .D(n814), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[14][27] ), .QN(n3446) );
  DFFARX1 \regfile_reg[15][27]  ( .D(n813), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[15][27] ), .QN(n3198) );
  DFFARX1 \regfile_reg[0][26]  ( .D(n812), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][26] ), .QN(n3066) );
  DFFARX1 \regfile_reg[1][26]  ( .D(n811), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][26] ), .QN(n3325) );
  DFFARX1 \regfile_reg[2][26]  ( .D(n810), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[2][26] ), .QN(n3445) );
  DFFARX1 \regfile_reg[3][26]  ( .D(n809), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[3][26] ), .QN(n3197) );
  DFFARX1 \regfile_reg[4][26]  ( .D(n808), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[4][26] ), .QN(n3065) );
  DFFARX1 \regfile_reg[5][26]  ( .D(n807), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[5][26] ), .QN(n3324) );
  DFFARX1 \regfile_reg[6][26]  ( .D(n806), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[6][26] ), .QN(n3444) );
  DFFARX1 \regfile_reg[7][26]  ( .D(n805), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[7][26] ), .QN(n3196) );
  DFFARX1 \regfile_reg[8][26]  ( .D(n804), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[8][26] ), .QN(n3064) );
  DFFARX1 \regfile_reg[9][26]  ( .D(n803), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[9][26] ), .QN(n3323) );
  DFFARX1 \regfile_reg[10][26]  ( .D(n802), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[10][26] ), .QN(n3443) );
  DFFARX1 \regfile_reg[11][26]  ( .D(n801), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[11][26] ), .QN(n3195) );
  DFFARX1 \regfile_reg[12][26]  ( .D(n800), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[12][26] ), .QN(n3063) );
  DFFARX1 \regfile_reg[13][26]  ( .D(n799), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[13][26] ), .QN(n3322) );
  DFFARX1 \regfile_reg[14][26]  ( .D(n798), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[14][26] ), .QN(n3442) );
  DFFARX1 \regfile_reg[15][26]  ( .D(n797), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[15][26] ), .QN(n3194) );
  DFFARX1 \regfile_reg[0][25]  ( .D(n796), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[0][25] ), .QN(n3062) );
  DFFARX1 \regfile_reg[1][25]  ( .D(n795), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[1][25] ), .QN(n3321) );
  DFFARX1 \regfile_reg[2][25]  ( .D(n794), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[2][25] ), .QN(n3441) );
  DFFARX1 \regfile_reg[3][25]  ( .D(n793), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[3][25] ), .QN(n3193) );
  DFFARX1 \regfile_reg[4][25]  ( .D(n792), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][25] ), .QN(n3061) );
  DFFARX1 \regfile_reg[5][25]  ( .D(n791), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][25] ), .QN(n3320) );
  DFFARX1 \regfile_reg[6][25]  ( .D(n790), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[6][25] ), .QN(n3440) );
  DFFARX1 \regfile_reg[7][25]  ( .D(n789), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][25] ), .QN(n3192) );
  DFFARX1 \regfile_reg[8][25]  ( .D(n788), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][25] ), .QN(n3060) );
  DFFARX1 \regfile_reg[9][25]  ( .D(n787), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[9][25] ), .QN(n3319) );
  DFFARX1 \regfile_reg[10][25]  ( .D(n786), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[10][25] ), .QN(n3439) );
  DFFARX1 \regfile_reg[11][25]  ( .D(n785), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[11][25] ), .QN(n3191) );
  DFFARX1 \regfile_reg[12][25]  ( .D(n784), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[12][25] ), .QN(n3059) );
  DFFARX1 \regfile_reg[13][25]  ( .D(n783), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[13][25] ), .QN(n3318) );
  DFFARX1 \regfile_reg[14][25]  ( .D(n782), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[14][25] ), .QN(n3438) );
  DFFARX1 \regfile_reg[15][25]  ( .D(n781), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[15][25] ), .QN(n3190) );
  DFFARX1 \regfile_reg[0][24]  ( .D(n780), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][24] ), .QN(n3058) );
  DFFARX1 \regfile_reg[1][24]  ( .D(n779), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][24] ), .QN(n3317) );
  DFFARX1 \regfile_reg[2][24]  ( .D(n778), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[2][24] ), .QN(n3437) );
  DFFARX1 \regfile_reg[3][24]  ( .D(n777), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[3][24] ), .QN(n3189) );
  DFFARX1 \regfile_reg[4][24]  ( .D(n776), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[4][24] ), .QN(n3057) );
  DFFARX1 \regfile_reg[5][24]  ( .D(n775), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[5][24] ), .QN(n3316) );
  DFFARX1 \regfile_reg[6][24]  ( .D(n774), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[6][24] ), .QN(n3436) );
  DFFARX1 \regfile_reg[7][24]  ( .D(n773), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[7][24] ), .QN(n3188) );
  DFFARX1 \regfile_reg[8][24]  ( .D(n772), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][24] ), .QN(n3056) );
  DFFARX1 \regfile_reg[9][24]  ( .D(n771), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[9][24] ), .QN(n3315) );
  DFFARX1 \regfile_reg[10][24]  ( .D(n770), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[10][24] ), .QN(n3435) );
  DFFARX1 \regfile_reg[11][24]  ( .D(n769), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[11][24] ), .QN(n3187) );
  DFFARX1 \regfile_reg[12][24]  ( .D(n768), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[12][24] ), .QN(n3055) );
  DFFARX1 \regfile_reg[13][24]  ( .D(n767), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][24] ), .QN(n3314) );
  DFFARX1 \regfile_reg[14][24]  ( .D(n766), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[14][24] ), .QN(n3434) );
  DFFARX1 \regfile_reg[15][24]  ( .D(n765), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[15][24] ), .QN(n3186) );
  DFFARX1 \regfile_reg[0][23]  ( .D(n764), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[0][23] ), .QN(n3054) );
  DFFARX1 \regfile_reg[1][23]  ( .D(n763), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[1][23] ), .QN(n3313) );
  DFFARX1 \regfile_reg[2][23]  ( .D(n762), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[2][23] ), .QN(n3433) );
  DFFARX1 \regfile_reg[3][23]  ( .D(n761), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[3][23] ), .QN(n3185) );
  DFFARX1 \regfile_reg[4][23]  ( .D(n760), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][23] ), .QN(n3053) );
  DFFARX1 \regfile_reg[5][23]  ( .D(n759), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][23] ), .QN(n3312) );
  DFFARX1 \regfile_reg[6][23]  ( .D(n758), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[6][23] ), .QN(n3432) );
  DFFARX1 \regfile_reg[7][23]  ( .D(n757), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][23] ), .QN(n3184) );
  DFFARX1 \regfile_reg[8][23]  ( .D(n756), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][23] ), .QN(n3052) );
  DFFARX1 \regfile_reg[9][23]  ( .D(n755), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[9][23] ), .QN(n3311) );
  DFFARX1 \regfile_reg[10][23]  ( .D(n754), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[10][23] ), .QN(n3431) );
  DFFARX1 \regfile_reg[11][23]  ( .D(n753), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[11][23] ), .QN(n3183) );
  DFFARX1 \regfile_reg[12][23]  ( .D(n752), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[12][23] ), .QN(n3051) );
  DFFARX1 \regfile_reg[13][23]  ( .D(n751), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[13][23] ), .QN(n3310) );
  DFFARX1 \regfile_reg[14][23]  ( .D(n750), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[14][23] ), .QN(n3430) );
  DFFARX1 \regfile_reg[15][23]  ( .D(n749), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[15][23] ), .QN(n3182) );
  DFFARX1 \regfile_reg[0][22]  ( .D(n748), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[0][22] ), .QN(n3050) );
  DFFARX1 \regfile_reg[1][22]  ( .D(n747), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][22] ), .QN(n3309) );
  DFFARX1 \regfile_reg[2][22]  ( .D(n746), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[2][22] ), .QN(n3429) );
  DFFARX1 \regfile_reg[3][22]  ( .D(n745), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[3][22] ), .QN(n3181) );
  DFFARX1 \regfile_reg[4][22]  ( .D(n744), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[4][22] ), .QN(n3049) );
  DFFARX1 \regfile_reg[5][22]  ( .D(n743), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[5][22] ), .QN(n3308) );
  DFFARX1 \regfile_reg[6][22]  ( .D(n742), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[6][22] ), .QN(n3428) );
  DFFARX1 \regfile_reg[7][22]  ( .D(n741), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[7][22] ), .QN(n3180) );
  DFFARX1 \regfile_reg[8][22]  ( .D(n740), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][22] ), .QN(n3048) );
  DFFARX1 \regfile_reg[9][22]  ( .D(n739), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[9][22] ), .QN(n3307) );
  DFFARX1 \regfile_reg[10][22]  ( .D(n738), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[10][22] ), .QN(n3427) );
  DFFARX1 \regfile_reg[11][22]  ( .D(n737), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[11][22] ), .QN(n3179) );
  DFFARX1 \regfile_reg[12][22]  ( .D(n736), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[12][22] ), .QN(n3047) );
  DFFARX1 \regfile_reg[13][22]  ( .D(n735), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][22] ), .QN(n3306) );
  DFFARX1 \regfile_reg[14][22]  ( .D(n734), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[14][22] ), .QN(n3426) );
  DFFARX1 \regfile_reg[15][22]  ( .D(n733), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[15][22] ), .QN(n3178) );
  DFFARX1 \regfile_reg[0][21]  ( .D(n732), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[0][21] ), .QN(n3046) );
  DFFARX1 \regfile_reg[1][21]  ( .D(n731), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[1][21] ), .QN(n3305) );
  DFFARX1 \regfile_reg[2][21]  ( .D(n730), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[2][21] ), .QN(n3425) );
  DFFARX1 \regfile_reg[3][21]  ( .D(n729), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[3][21] ), .QN(n3177) );
  DFFARX1 \regfile_reg[4][21]  ( .D(n728), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][21] ), .QN(n3045) );
  DFFARX1 \regfile_reg[5][21]  ( .D(n727), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][21] ), .QN(n3304) );
  DFFARX1 \regfile_reg[6][21]  ( .D(n726), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[6][21] ), .QN(n3424) );
  DFFARX1 \regfile_reg[7][21]  ( .D(n725), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][21] ), .QN(n3176) );
  DFFARX1 \regfile_reg[8][21]  ( .D(n724), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][21] ), .QN(n3044) );
  DFFARX1 \regfile_reg[9][21]  ( .D(n723), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[9][21] ), .QN(n3303) );
  DFFARX1 \regfile_reg[10][21]  ( .D(n722), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[10][21] ), .QN(n3423) );
  DFFARX1 \regfile_reg[11][21]  ( .D(n721), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[11][21] ), .QN(n3175) );
  DFFARX1 \regfile_reg[12][21]  ( .D(n720), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[12][21] ), .QN(n3043) );
  DFFARX1 \regfile_reg[13][21]  ( .D(n719), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[13][21] ), .QN(n3302) );
  DFFARX1 \regfile_reg[14][21]  ( .D(n718), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[14][21] ), .QN(n3422) );
  DFFARX1 \regfile_reg[15][21]  ( .D(n717), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[15][21] ), .QN(n3174) );
  DFFARX1 \regfile_reg[0][20]  ( .D(n716), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[0][20] ), .QN(n3042) );
  DFFARX1 \regfile_reg[1][20]  ( .D(n715), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][20] ), .QN(n3301) );
  DFFARX1 \regfile_reg[2][20]  ( .D(n714), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[2][20] ), .QN(n3421) );
  DFFARX1 \regfile_reg[3][20]  ( .D(n713), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[3][20] ), .QN(n3173) );
  DFFARX1 \regfile_reg[4][20]  ( .D(n712), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[4][20] ), .QN(n3041) );
  DFFARX1 \regfile_reg[5][20]  ( .D(n711), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[5][20] ), .QN(n3300) );
  DFFARX1 \regfile_reg[6][20]  ( .D(n710), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[6][20] ), .QN(n3420) );
  DFFARX1 \regfile_reg[7][20]  ( .D(n709), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[7][20] ), .QN(n3172) );
  DFFARX1 \regfile_reg[8][20]  ( .D(n708), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][20] ), .QN(n3040) );
  DFFARX1 \regfile_reg[9][20]  ( .D(n707), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[9][20] ), .QN(n3299) );
  DFFARX1 \regfile_reg[10][20]  ( .D(n706), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[10][20] ), .QN(n3419) );
  DFFARX1 \regfile_reg[11][20]  ( .D(n705), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[11][20] ), .QN(n3171) );
  DFFARX1 \regfile_reg[12][20]  ( .D(n704), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[12][20] ), .QN(n3039) );
  DFFARX1 \regfile_reg[13][20]  ( .D(n703), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][20] ), .QN(n3298) );
  DFFARX1 \regfile_reg[14][20]  ( .D(n702), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[14][20] ), .QN(n3418) );
  DFFARX1 \regfile_reg[15][20]  ( .D(n701), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[15][20] ), .QN(n3170) );
  DFFARX1 \regfile_reg[0][19]  ( .D(n700), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[0][19] ), .QN(n3038) );
  DFFARX1 \regfile_reg[1][19]  ( .D(n699), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][19] ), .QN(n3297) );
  DFFARX1 \regfile_reg[2][19]  ( .D(n698), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[2][19] ), .QN(n3417) );
  DFFARX1 \regfile_reg[3][19]  ( .D(n697), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[3][19] ), .QN(n3169) );
  DFFARX1 \regfile_reg[4][19]  ( .D(n696), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[4][19] ), .QN(n3037) );
  DFFARX1 \regfile_reg[5][19]  ( .D(n695), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[5][19] ), .QN(n3296) );
  DFFARX1 \regfile_reg[6][19]  ( .D(n694), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[6][19] ), .QN(n3416) );
  DFFARX1 \regfile_reg[7][19]  ( .D(n693), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[7][19] ), .QN(n3168) );
  DFFARX1 \regfile_reg[8][19]  ( .D(n692), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][19] ), .QN(n3036) );
  DFFARX1 \regfile_reg[9][19]  ( .D(n691), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[9][19] ), .QN(n3295) );
  DFFARX1 \regfile_reg[10][19]  ( .D(n690), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[10][19] ), .QN(n3415) );
  DFFARX1 \regfile_reg[11][19]  ( .D(n689), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[11][19] ), .QN(n3167) );
  DFFARX1 \regfile_reg[12][19]  ( .D(n688), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[12][19] ), .QN(n3035) );
  DFFARX1 \regfile_reg[13][19]  ( .D(n687), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][19] ), .QN(n3294) );
  DFFARX1 \regfile_reg[14][19]  ( .D(n686), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[14][19] ), .QN(n3414) );
  DFFARX1 \regfile_reg[15][19]  ( .D(n685), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[15][19] ), .QN(n3166) );
  DFFARX1 \regfile_reg[0][18]  ( .D(n684), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[0][18] ), .QN(n3034) );
  DFFARX1 \regfile_reg[1][18]  ( .D(n683), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[1][18] ), .QN(n3293) );
  DFFARX1 \regfile_reg[2][18]  ( .D(n682), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[2][18] ), .QN(n3413) );
  DFFARX1 \regfile_reg[3][18]  ( .D(n681), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[3][18] ), .QN(n3165) );
  DFFARX1 \regfile_reg[4][18]  ( .D(n680), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][18] ), .QN(n3033) );
  DFFARX1 \regfile_reg[5][18]  ( .D(n679), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][18] ), .QN(n3292) );
  DFFARX1 \regfile_reg[6][18]  ( .D(n678), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[6][18] ), .QN(n3412) );
  DFFARX1 \regfile_reg[7][18]  ( .D(n677), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][18] ), .QN(n3164) );
  DFFARX1 \regfile_reg[8][18]  ( .D(n676), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][18] ), .QN(n3032) );
  DFFARX1 \regfile_reg[9][18]  ( .D(n675), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[9][18] ), .QN(n3291) );
  DFFARX1 \regfile_reg[10][18]  ( .D(n674), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[10][18] ), .QN(n3411) );
  DFFARX1 \regfile_reg[11][18]  ( .D(n673), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[11][18] ), .QN(n3163) );
  DFFARX1 \regfile_reg[12][18]  ( .D(n672), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[12][18] ), .QN(n3031) );
  DFFARX1 \regfile_reg[13][18]  ( .D(n671), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[13][18] ), .QN(n3290) );
  DFFARX1 \regfile_reg[14][18]  ( .D(n670), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[14][18] ), .QN(n3410) );
  DFFARX1 \regfile_reg[15][18]  ( .D(n669), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[15][18] ), .QN(n3162) );
  DFFARX1 \regfile_reg[0][17]  ( .D(n668), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[0][17] ), .QN(n3030) );
  DFFARX1 \regfile_reg[1][17]  ( .D(n667), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][17] ), .QN(n3289) );
  DFFARX1 \regfile_reg[2][17]  ( .D(n666), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[2][17] ), .QN(n3409) );
  DFFARX1 \regfile_reg[3][17]  ( .D(n665), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[3][17] ), .QN(n3161) );
  DFFARX1 \regfile_reg[4][17]  ( .D(n664), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[4][17] ), .QN(n3029) );
  DFFARX1 \regfile_reg[5][17]  ( .D(n663), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[5][17] ), .QN(n3288) );
  DFFARX1 \regfile_reg[6][17]  ( .D(n662), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[6][17] ), .QN(n3408) );
  DFFARX1 \regfile_reg[7][17]  ( .D(n661), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[7][17] ), .QN(n3160) );
  DFFARX1 \regfile_reg[8][17]  ( .D(n660), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][17] ), .QN(n3028) );
  DFFARX1 \regfile_reg[9][17]  ( .D(n659), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[9][17] ), .QN(n3287) );
  DFFARX1 \regfile_reg[10][17]  ( .D(n658), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[10][17] ), .QN(n3407) );
  DFFARX1 \regfile_reg[11][17]  ( .D(n657), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[11][17] ), .QN(n3159) );
  DFFARX1 \regfile_reg[12][17]  ( .D(n656), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[12][17] ), .QN(n3027) );
  DFFARX1 \regfile_reg[13][17]  ( .D(n655), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][17] ), .QN(n3286) );
  DFFARX1 \regfile_reg[14][17]  ( .D(n654), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[14][17] ), .QN(n3406) );
  DFFARX1 \regfile_reg[15][17]  ( .D(n653), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[15][17] ), .QN(n3158) );
  DFFARX1 \regfile_reg[0][16]  ( .D(n652), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][16] ), .QN(n3026) );
  DFFARX1 \regfile_reg[1][16]  ( .D(n651), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[1][16] ), .QN(n3285) );
  DFFARX1 \regfile_reg[2][16]  ( .D(n650), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[2][16] ), .QN(n3405) );
  DFFARX1 \regfile_reg[3][16]  ( .D(n649), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[3][16] ), .QN(n3157) );
  DFFARX1 \regfile_reg[4][16]  ( .D(n648), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][16] ), .QN(n3025) );
  DFFARX1 \regfile_reg[5][16]  ( .D(n647), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][16] ), .QN(n3284) );
  DFFARX1 \regfile_reg[6][16]  ( .D(n646), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[6][16] ), .QN(n3404) );
  DFFARX1 \regfile_reg[7][16]  ( .D(n645), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[7][16] ), .QN(n3156) );
  DFFARX1 \regfile_reg[8][16]  ( .D(n644), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][16] ), .QN(n3024) );
  DFFARX1 \regfile_reg[9][16]  ( .D(n643), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[9][16] ), .QN(n3283) );
  DFFARX1 \regfile_reg[10][16]  ( .D(n642), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[10][16] ), .QN(n3403) );
  DFFARX1 \regfile_reg[11][16]  ( .D(n641), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[11][16] ), .QN(n3155) );
  DFFARX1 \regfile_reg[12][16]  ( .D(n640), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[12][16] ), .QN(n3023) );
  DFFARX1 \regfile_reg[13][16]  ( .D(n639), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[13][16] ), .QN(n3282) );
  DFFARX1 \regfile_reg[14][16]  ( .D(n638), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[14][16] ), .QN(n3402) );
  DFFARX1 \regfile_reg[15][16]  ( .D(n637), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[15][16] ), .QN(n3154) );
  DFFARX1 \regfile_reg[0][15]  ( .D(n636), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[0][15] ), .QN(n3022) );
  DFFARX1 \regfile_reg[1][15]  ( .D(n635), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][15] ), .QN(n3281) );
  DFFARX1 \regfile_reg[2][15]  ( .D(n634), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[2][15] ), .QN(n3401) );
  DFFARX1 \regfile_reg[3][15]  ( .D(n633), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[3][15] ), .QN(n3153) );
  DFFARX1 \regfile_reg[4][15]  ( .D(n632), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[4][15] ), .QN(n3021) );
  DFFARX1 \regfile_reg[5][15]  ( .D(n631), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[5][15] ), .QN(n3280) );
  DFFARX1 \regfile_reg[6][15]  ( .D(n630), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[6][15] ), .QN(n3400) );
  DFFARX1 \regfile_reg[7][15]  ( .D(n629), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[7][15] ), .QN(n3152) );
  DFFARX1 \regfile_reg[8][15]  ( .D(n628), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][15] ), .QN(n3020) );
  DFFARX1 \regfile_reg[9][15]  ( .D(n627), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[9][15] ), .QN(n3279) );
  DFFARX1 \regfile_reg[10][15]  ( .D(n626), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[10][15] ), .QN(n3399) );
  DFFARX1 \regfile_reg[11][15]  ( .D(n625), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[11][15] ), .QN(n3151) );
  DFFARX1 \regfile_reg[12][15]  ( .D(n624), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[12][15] ), .QN(n3019) );
  DFFARX1 \regfile_reg[13][15]  ( .D(n623), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][15] ), .QN(n3278) );
  DFFARX1 \regfile_reg[14][15]  ( .D(n622), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[14][15] ), .QN(n3398) );
  DFFARX1 \regfile_reg[15][15]  ( .D(n621), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[15][15] ), .QN(n3150) );
  DFFARX1 \regfile_reg[0][14]  ( .D(n620), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][14] ), .QN(n3018) );
  DFFARX1 \regfile_reg[1][14]  ( .D(n619), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[1][14] ), .QN(n3277) );
  DFFARX1 \regfile_reg[2][14]  ( .D(n618), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[2][14] ), .QN(n3397) );
  DFFARX1 \regfile_reg[3][14]  ( .D(n617), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[3][14] ), .QN(n3149) );
  DFFARX1 \regfile_reg[4][14]  ( .D(n616), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[4][14] ), .QN(n3017) );
  DFFARX1 \regfile_reg[5][14]  ( .D(n615), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][14] ), .QN(n3276) );
  DFFARX1 \regfile_reg[6][14]  ( .D(n614), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[6][14] ), .QN(n3396) );
  DFFARX1 \regfile_reg[7][14]  ( .D(n613), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[7][14] ), .QN(n3148) );
  DFFARX1 \regfile_reg[8][14]  ( .D(n612), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][14] ), .QN(n3016) );
  DFFARX1 \regfile_reg[9][14]  ( .D(n611), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[9][14] ), .QN(n3275) );
  DFFARX1 \regfile_reg[10][14]  ( .D(n610), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[10][14] ), .QN(n3395) );
  DFFARX1 \regfile_reg[11][14]  ( .D(n609), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[11][14] ), .QN(n3147) );
  DFFARX1 \regfile_reg[12][14]  ( .D(n608), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[12][14] ), .QN(n3015) );
  DFFARX1 \regfile_reg[13][14]  ( .D(n607), .CLK(clk), .RSTB(n3748), .Q(
        \regfile[13][14] ), .QN(n3274) );
  DFFARX1 \regfile_reg[14][14]  ( .D(n606), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[14][14] ), .QN(n3394) );
  DFFARX1 \regfile_reg[15][14]  ( .D(n605), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[15][14] ), .QN(n3146) );
  DFFARX1 \regfile_reg[0][13]  ( .D(n604), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][13] ), .QN(n3014) );
  DFFARX1 \regfile_reg[1][13]  ( .D(n603), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][13] ), .QN(n3273) );
  DFFARX1 \regfile_reg[2][13]  ( .D(n602), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[2][13] ), .QN(n3393) );
  DFFARX1 \regfile_reg[3][13]  ( .D(n601), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[3][13] ), .QN(n3145) );
  DFFARX1 \regfile_reg[4][13]  ( .D(n600), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[4][13] ), .QN(n3013) );
  DFFARX1 \regfile_reg[5][13]  ( .D(n599), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[5][13] ), .QN(n3272) );
  DFFARX1 \regfile_reg[6][13]  ( .D(n598), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[6][13] ), .QN(n3392) );
  DFFARX1 \regfile_reg[7][13]  ( .D(n597), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[7][13] ), .QN(n3144) );
  DFFARX1 \regfile_reg[8][13]  ( .D(n596), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][13] ), .QN(n3012) );
  DFFARX1 \regfile_reg[9][13]  ( .D(n595), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[9][13] ), .QN(n3271) );
  DFFARX1 \regfile_reg[10][13]  ( .D(n594), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[10][13] ), .QN(n3391) );
  DFFARX1 \regfile_reg[11][13]  ( .D(n593), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[11][13] ), .QN(n3143) );
  DFFARX1 \regfile_reg[12][13]  ( .D(n592), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[12][13] ), .QN(n3011) );
  DFFARX1 \regfile_reg[13][13]  ( .D(n591), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][13] ), .QN(n3270) );
  DFFARX1 \regfile_reg[14][13]  ( .D(n590), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[14][13] ), .QN(n3390) );
  DFFARX1 \regfile_reg[15][13]  ( .D(n589), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[15][13] ), .QN(n3142) );
  DFFARX1 \regfile_reg[0][12]  ( .D(n588), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][12] ), .QN(n3010) );
  DFFARX1 \regfile_reg[1][12]  ( .D(n587), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[1][12] ), .QN(n3269) );
  DFFARX1 \regfile_reg[2][12]  ( .D(n586), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[2][12] ), .QN(n3389) );
  DFFARX1 \regfile_reg[3][12]  ( .D(n585), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[3][12] ), .QN(n3141) );
  DFFARX1 \regfile_reg[4][12]  ( .D(n584), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[4][12] ), .QN(n3009) );
  DFFARX1 \regfile_reg[5][12]  ( .D(n583), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][12] ), .QN(n3268) );
  DFFARX1 \regfile_reg[6][12]  ( .D(n582), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[6][12] ), .QN(n3388) );
  DFFARX1 \regfile_reg[7][12]  ( .D(n581), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[7][12] ), .QN(n3140) );
  DFFARX1 \regfile_reg[8][12]  ( .D(n580), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][12] ), .QN(n3008) );
  DFFARX1 \regfile_reg[9][12]  ( .D(n579), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[9][12] ), .QN(n3267) );
  DFFARX1 \regfile_reg[10][12]  ( .D(n578), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[10][12] ), .QN(n3387) );
  DFFARX1 \regfile_reg[11][12]  ( .D(n577), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[11][12] ), .QN(n3139) );
  DFFARX1 \regfile_reg[12][12]  ( .D(n576), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[12][12] ), .QN(n3007) );
  DFFARX1 \regfile_reg[13][12]  ( .D(n575), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[13][12] ), .QN(n3266) );
  DFFARX1 \regfile_reg[14][12]  ( .D(n574), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[14][12] ), .QN(n3386) );
  DFFARX1 \regfile_reg[15][12]  ( .D(n573), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[15][12] ), .QN(n3138) );
  DFFARX1 \regfile_reg[0][11]  ( .D(n572), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][11] ), .QN(n3006) );
  DFFARX1 \regfile_reg[1][11]  ( .D(n571), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][11] ), .QN(n3265) );
  DFFARX1 \regfile_reg[2][11]  ( .D(n570), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[2][11] ), .QN(n3385) );
  DFFARX1 \regfile_reg[3][11]  ( .D(n569), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[3][11] ), .QN(n3137) );
  DFFARX1 \regfile_reg[4][11]  ( .D(n568), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[4][11] ), .QN(n3005) );
  DFFARX1 \regfile_reg[5][11]  ( .D(n567), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[5][11] ), .QN(n3264) );
  DFFARX1 \regfile_reg[6][11]  ( .D(n566), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[6][11] ), .QN(n3384) );
  DFFARX1 \regfile_reg[7][11]  ( .D(n565), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[7][11] ), .QN(n3136) );
  DFFARX1 \regfile_reg[8][11]  ( .D(n564), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[8][11] ), .QN(n3004) );
  DFFARX1 \regfile_reg[9][11]  ( .D(n563), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[9][11] ), .QN(n3263) );
  DFFARX1 \regfile_reg[10][11]  ( .D(n562), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[10][11] ), .QN(n3383) );
  DFFARX1 \regfile_reg[11][11]  ( .D(n561), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[11][11] ), .QN(n3135) );
  DFFARX1 \regfile_reg[12][11]  ( .D(n560), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[12][11] ), .QN(n3003) );
  DFFARX1 \regfile_reg[13][11]  ( .D(n559), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[13][11] ), .QN(n3262) );
  DFFARX1 \regfile_reg[14][11]  ( .D(n558), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[14][11] ), .QN(n3382) );
  DFFARX1 \regfile_reg[15][11]  ( .D(n557), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[15][11] ), .QN(n3134) );
  DFFARX1 \regfile_reg[0][10]  ( .D(n556), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][10] ), .QN(n3002) );
  DFFARX1 \regfile_reg[1][10]  ( .D(n555), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[1][10] ), .QN(n3261) );
  DFFARX1 \regfile_reg[2][10]  ( .D(n554), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[2][10] ), .QN(n3381) );
  DFFARX1 \regfile_reg[3][10]  ( .D(n553), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[3][10] ), .QN(n3133) );
  DFFARX1 \regfile_reg[4][10]  ( .D(n552), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[4][10] ), .QN(n3001) );
  DFFARX1 \regfile_reg[5][10]  ( .D(n551), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[5][10] ), .QN(n3260) );
  DFFARX1 \regfile_reg[6][10]  ( .D(n550), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[6][10] ), .QN(n3380) );
  DFFARX1 \regfile_reg[7][10]  ( .D(n549), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[7][10] ), .QN(n3132) );
  DFFARX1 \regfile_reg[8][10]  ( .D(n548), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[8][10] ), .QN(n3000) );
  DFFARX1 \regfile_reg[9][10]  ( .D(n547), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[9][10] ), .QN(n3259) );
  DFFARX1 \regfile_reg[10][10]  ( .D(n546), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[10][10] ), .QN(n3379) );
  DFFARX1 \regfile_reg[11][10]  ( .D(n545), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[11][10] ), .QN(n3131) );
  DFFARX1 \regfile_reg[12][10]  ( .D(n544), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[12][10] ), .QN(n2999) );
  DFFARX1 \regfile_reg[13][10]  ( .D(n543), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[13][10] ), .QN(n3258) );
  DFFARX1 \regfile_reg[14][10]  ( .D(n542), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[14][10] ), .QN(n3378) );
  DFFARX1 \regfile_reg[15][10]  ( .D(n541), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[15][10] ), .QN(n3130) );
  DFFARX1 \regfile_reg[0][9]  ( .D(n540), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[0][9] ), .QN(n2998) );
  DFFARX1 \regfile_reg[1][9]  ( .D(n539), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[1][9] ), .QN(n3257) );
  DFFARX1 \regfile_reg[2][9]  ( .D(n538), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[2][9] ), .QN(n3377) );
  DFFARX1 \regfile_reg[3][9]  ( .D(n537), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[3][9] ), .QN(n3129) );
  DFFARX1 \regfile_reg[4][9]  ( .D(n536), .CLK(clk), .RSTB(n3742), .Q(
        \regfile[4][9] ), .QN(n2997) );
  DFFARX1 \regfile_reg[5][9]  ( .D(n535), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[5][9] ), .QN(n3256) );
  DFFARX1 \regfile_reg[6][9]  ( .D(n534), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[6][9] ), .QN(n3376) );
  DFFARX1 \regfile_reg[7][9]  ( .D(n533), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][9] ), .QN(n3128) );
  DFFARX1 \regfile_reg[8][9]  ( .D(n532), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[8][9] ), .QN(n2996) );
  DFFARX1 \regfile_reg[9][9]  ( .D(n531), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[9][9] ), .QN(n3255) );
  DFFARX1 \regfile_reg[10][9]  ( .D(n530), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[10][9] ), .QN(n3375) );
  DFFARX1 \regfile_reg[11][9]  ( .D(n529), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[11][9] ), .QN(n3127) );
  DFFARX1 \regfile_reg[12][9]  ( .D(n528), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[12][9] ), .QN(n2995) );
  DFFARX1 \regfile_reg[13][9]  ( .D(n527), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[13][9] ), .QN(n3254) );
  DFFARX1 \regfile_reg[14][9]  ( .D(n526), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[14][9] ), .QN(n3374) );
  DFFARX1 \regfile_reg[15][9]  ( .D(n525), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[15][9] ), .QN(n3126) );
  DFFARX1 \regfile_reg[0][8]  ( .D(n524), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[0][8] ), .QN(n2994) );
  DFFARX1 \regfile_reg[1][8]  ( .D(n523), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[1][8] ), .QN(n3253) );
  DFFARX1 \regfile_reg[2][8]  ( .D(n522), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[2][8] ), .QN(n3373) );
  DFFARX1 \regfile_reg[3][8]  ( .D(n521), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[3][8] ), .QN(n3125) );
  DFFARX1 \regfile_reg[4][8]  ( .D(n520), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[4][8] ), .QN(n2993) );
  DFFARX1 \regfile_reg[5][8]  ( .D(n519), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[5][8] ), .QN(n3252) );
  DFFARX1 \regfile_reg[6][8]  ( .D(n518), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[6][8] ), .QN(n3372) );
  DFFARX1 \regfile_reg[7][8]  ( .D(n517), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[7][8] ), .QN(n3124) );
  DFFARX1 \regfile_reg[8][8]  ( .D(n516), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[8][8] ), .QN(n2992) );
  DFFARX1 \regfile_reg[9][8]  ( .D(n515), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[9][8] ), .QN(n3251) );
  DFFARX1 \regfile_reg[10][8]  ( .D(n514), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[10][8] ), .QN(n3371) );
  DFFARX1 \regfile_reg[11][8]  ( .D(n513), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[11][8] ), .QN(n3123) );
  DFFARX1 \regfile_reg[12][8]  ( .D(n512), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[12][8] ), .QN(n2991) );
  DFFARX1 \regfile_reg[13][8]  ( .D(n511), .CLK(clk), .RSTB(n3763), .Q(
        \regfile[13][8] ), .QN(n3250) );
  DFFARX1 \regfile_reg[14][8]  ( .D(n510), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[14][8] ), .QN(n3370) );
  DFFARX1 \regfile_reg[15][8]  ( .D(n509), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[15][8] ), .QN(n3122) );
  DFFARX1 \regfile_reg[0][7]  ( .D(n508), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[0][7] ), .QN(n2990) );
  DFFARX1 \regfile_reg[1][7]  ( .D(n507), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[1][7] ), .QN(n3249) );
  DFFARX1 \regfile_reg[2][7]  ( .D(n506), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[2][7] ), .QN(n3369) );
  DFFARX1 \regfile_reg[3][7]  ( .D(n505), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[3][7] ), .QN(n3121) );
  DFFARX1 \regfile_reg[4][7]  ( .D(n504), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][7] ), .QN(n2989) );
  DFFARX1 \regfile_reg[5][7]  ( .D(n503), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[5][7] ), .QN(n3248) );
  DFFARX1 \regfile_reg[6][7]  ( .D(n502), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[6][7] ), .QN(n3368) );
  DFFARX1 \regfile_reg[7][7]  ( .D(n501), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][7] ), .QN(n3120) );
  DFFARX1 \regfile_reg[8][7]  ( .D(n500), .CLK(clk), .RSTB(n3737), .Q(
        \regfile[8][7] ), .QN(n2988) );
  DFFARX1 \regfile_reg[9][7]  ( .D(n499), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[9][7] ), .QN(n3247) );
  DFFARX1 \regfile_reg[10][7]  ( .D(n498), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[10][7] ), .QN(n3367) );
  DFFARX1 \regfile_reg[11][7]  ( .D(n497), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[11][7] ), .QN(n3119) );
  DFFARX1 \regfile_reg[12][7]  ( .D(n496), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[12][7] ), .QN(n2987) );
  DFFARX1 \regfile_reg[13][7]  ( .D(n495), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[13][7] ), .QN(n3246) );
  DFFARX1 \regfile_reg[14][7]  ( .D(n494), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[14][7] ), .QN(n3366) );
  DFFARX1 \regfile_reg[15][7]  ( .D(n493), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[15][7] ), .QN(n3118) );
  DFFARX1 \regfile_reg[0][6]  ( .D(n492), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[0][6] ), .QN(n2986) );
  DFFARX1 \regfile_reg[1][6]  ( .D(n491), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[1][6] ), .QN(n3245) );
  DFFARX1 \regfile_reg[2][6]  ( .D(n490), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[2][6] ), .QN(n3365) );
  DFFARX1 \regfile_reg[3][6]  ( .D(n489), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[3][6] ), .QN(n3117) );
  DFFARX1 \regfile_reg[4][6]  ( .D(n488), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[4][6] ), .QN(n2985) );
  DFFARX1 \regfile_reg[5][6]  ( .D(n487), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[5][6] ), .QN(n3244) );
  DFFARX1 \regfile_reg[6][6]  ( .D(n486), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[6][6] ), .QN(n3364) );
  DFFARX1 \regfile_reg[7][6]  ( .D(n485), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[7][6] ), .QN(n3116) );
  DFFARX1 \regfile_reg[8][6]  ( .D(n484), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[8][6] ), .QN(n2984) );
  DFFARX1 \regfile_reg[9][6]  ( .D(n483), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[9][6] ), .QN(n3243) );
  DFFARX1 \regfile_reg[10][6]  ( .D(n482), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[10][6] ), .QN(n3363) );
  DFFARX1 \regfile_reg[11][6]  ( .D(n481), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[11][6] ), .QN(n3115) );
  DFFARX1 \regfile_reg[12][6]  ( .D(n480), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[12][6] ), .QN(n2983) );
  DFFARX1 \regfile_reg[13][6]  ( .D(n479), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][6] ), .QN(n3242) );
  DFFARX1 \regfile_reg[14][6]  ( .D(n478), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[14][6] ), .QN(n3362) );
  DFFARX1 \regfile_reg[15][6]  ( .D(n477), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[15][6] ), .QN(n3114) );
  DFFARX1 \regfile_reg[0][5]  ( .D(n476), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[0][5] ), .QN(n2982) );
  DFFARX1 \regfile_reg[1][5]  ( .D(n475), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[1][5] ), .QN(n3241) );
  DFFARX1 \regfile_reg[2][5]  ( .D(n474), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[2][5] ), .QN(n3361) );
  DFFARX1 \regfile_reg[3][5]  ( .D(n473), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[3][5] ), .QN(n3113) );
  DFFARX1 \regfile_reg[4][5]  ( .D(n472), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][5] ), .QN(n2981) );
  DFFARX1 \regfile_reg[5][5]  ( .D(n471), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[5][5] ), .QN(n3240) );
  DFFARX1 \regfile_reg[6][5]  ( .D(n470), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[6][5] ), .QN(n3360) );
  DFFARX1 \regfile_reg[7][5]  ( .D(n469), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][5] ), .QN(n3112) );
  DFFARX1 \regfile_reg[8][5]  ( .D(n468), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][5] ), .QN(n2980) );
  DFFARX1 \regfile_reg[9][5]  ( .D(n467), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[9][5] ), .QN(n3239) );
  DFFARX1 \regfile_reg[10][5]  ( .D(n466), .CLK(clk), .RSTB(n3734), .Q(
        \regfile[10][5] ), .QN(n3359) );
  DFFARX1 \regfile_reg[11][5]  ( .D(n465), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[11][5] ), .QN(n3111) );
  DFFARX1 \regfile_reg[12][5]  ( .D(n464), .CLK(clk), .RSTB(n3736), .Q(
        \regfile[12][5] ), .QN(n2979) );
  DFFARX1 \regfile_reg[13][5]  ( .D(n463), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[13][5] ), .QN(n3238) );
  DFFARX1 \regfile_reg[14][5]  ( .D(n462), .CLK(clk), .RSTB(n3750), .Q(
        \regfile[14][5] ), .QN(n3358) );
  DFFARX1 \regfile_reg[15][5]  ( .D(n461), .CLK(clk), .RSTB(n3752), .Q(
        \regfile[15][5] ), .QN(n3110) );
  DFFARX1 \regfile_reg[0][4]  ( .D(n460), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[0][4] ), .QN(n2978) );
  DFFARX1 \regfile_reg[1][4]  ( .D(n459), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[1][4] ), .QN(n3237) );
  DFFARX1 \regfile_reg[2][4]  ( .D(n458), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[2][4] ), .QN(n3357) );
  DFFARX1 \regfile_reg[3][4]  ( .D(n457), .CLK(clk), .RSTB(n3725), .Q(
        \regfile[3][4] ), .QN(n3109) );
  DFFARX1 \regfile_reg[4][4]  ( .D(n456), .CLK(clk), .RSTB(n3726), .Q(
        \regfile[4][4] ), .QN(n2977) );
  DFFARX1 \regfile_reg[5][4]  ( .D(n455), .CLK(clk), .RSTB(n3728), .Q(
        \regfile[5][4] ), .QN(n3236) );
  DFFARX1 \regfile_reg[6][4]  ( .D(n454), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[6][4] ), .QN(n3356) );
  DFFARX1 \regfile_reg[7][4]  ( .D(n453), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[7][4] ), .QN(n3108) );
  DFFARX1 \regfile_reg[8][4]  ( .D(n452), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][4] ), .QN(n2976) );
  DFFARX1 \regfile_reg[9][4]  ( .D(n451), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[9][4] ), .QN(n3235) );
  DFFARX1 \regfile_reg[10][4]  ( .D(n450), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[10][4] ), .QN(n3355) );
  DFFARX1 \regfile_reg[11][4]  ( .D(n449), .CLK(clk), .RSTB(n3760), .Q(
        \regfile[11][4] ), .QN(n3107) );
  DFFARX1 \regfile_reg[12][4]  ( .D(n448), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[12][4] ), .QN(n2975) );
  DFFARX1 \regfile_reg[13][4]  ( .D(n447), .CLK(clk), .RSTB(n3762), .Q(
        \regfile[13][4] ), .QN(n3234) );
  DFFARX1 \regfile_reg[14][4]  ( .D(n446), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[14][4] ), .QN(n3221) );
  DFFASX1 \regfile_reg[15][4]  ( .D(n445), .CLK(clk), .SETB(n3765), .Q(
        \regfile[15][4] ), .QN(n3469) );
  DFFARX1 \regfile_reg[0][3]  ( .D(n444), .CLK(clk), .RSTB(n3735), .Q(
        \regfile[0][3] ), .QN(n2974) );
  DFFARX1 \regfile_reg[1][3]  ( .D(n443), .CLK(clk), .RSTB(n3753), .Q(
        \regfile[1][3] ), .QN(n3233) );
  DFFARX1 \regfile_reg[2][3]  ( .D(n442), .CLK(clk), .RSTB(n3754), .Q(
        \regfile[2][3] ), .QN(n3354) );
  DFFARX1 \regfile_reg[3][3]  ( .D(n441), .CLK(clk), .RSTB(n3744), .Q(
        \regfile[3][3] ), .QN(n3106) );
  DFFARX1 \regfile_reg[4][3]  ( .D(n440), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][3] ), .QN(n2973) );
  DFFARX1 \regfile_reg[5][3]  ( .D(n439), .CLK(clk), .RSTB(n3741), .Q(
        \regfile[5][3] ), .QN(n3232) );
  DFFARX1 \regfile_reg[6][3]  ( .D(n438), .CLK(clk), .RSTB(n3740), .Q(
        \regfile[6][3] ), .QN(n3220) );
  DFFASX1 \regfile_reg[7][3]  ( .D(n437), .CLK(clk), .SETB(n3764), .Q(
        \regfile[7][3] ), .QN(n3468) );
  DFFASX1 \regfile_reg[8][3]  ( .D(n436), .CLK(clk), .SETB(n3764), .Q(
        \regfile[8][3] ), .QN(n3094) );
  DFFASX1 \regfile_reg[9][3]  ( .D(n435), .CLK(clk), .SETB(n3764), .Q(
        \regfile[9][3] ), .QN(n3353) );
  DFFASX1 \regfile_reg[10][3]  ( .D(n434), .CLK(clk), .SETB(n3764), .Q(
        \regfile[10][3] ), .QN(n3481) );
  DFFASX1 \regfile_reg[11][3]  ( .D(n433), .CLK(clk), .SETB(n3764), .Q(
        \regfile[11][3] ), .QN(n3222) );
  DFFASX1 \regfile_reg[12][3]  ( .D(n432), .CLK(clk), .SETB(n3764), .Q(
        \regfile[12][3] ), .QN(n3093) );
  DFFASX1 \regfile_reg[13][3]  ( .D(n431), .CLK(clk), .SETB(n3764), .Q(
        \regfile[13][3] ), .QN(n3352) );
  DFFASX1 \regfile_reg[14][3]  ( .D(n430), .CLK(clk), .SETB(n3764), .Q(
        \regfile[14][3] ), .QN(n3480) );
  DFFARX1 \regfile_reg[15][3]  ( .D(n429), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[15][3] ), .QN(n3105) );
  DFFARX1 \regfile_reg[0][2]  ( .D(n428), .CLK(clk), .RSTB(n3757), .Q(
        \regfile[0][2] ), .QN(n2972) );
  DFFARX1 \regfile_reg[1][2]  ( .D(n427), .CLK(clk), .RSTB(n3747), .Q(
        \regfile[1][2] ), .QN(n3231) );
  DFFARX1 \regfile_reg[2][2]  ( .D(n426), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[2][2] ), .QN(n3219) );
  DFFASX1 \regfile_reg[3][2]  ( .D(n425), .CLK(clk), .SETB(n3764), .Q(
        \regfile[3][2] ), .QN(n3467) );
  DFFASX1 \regfile_reg[4][2]  ( .D(n424), .CLK(clk), .SETB(n3764), .Q(
        \regfile[4][2] ), .QN(n3092) );
  DFFASX1 \regfile_reg[5][2]  ( .D(n423), .CLK(clk), .SETB(n3764), .Q(
        \regfile[5][2] ), .QN(n3351) );
  DFFASX1 \regfile_reg[6][2]  ( .D(n422), .CLK(clk), .SETB(n3764), .Q(
        \regfile[6][2] ), .QN(n3479) );
  DFFARX1 \regfile_reg[7][2]  ( .D(n421), .CLK(clk), .RSTB(n3730), .Q(
        \regfile[7][2] ), .QN(n3104) );
  DFFARX1 \regfile_reg[8][2]  ( .D(n420), .CLK(clk), .RSTB(n3731), .Q(
        \regfile[8][2] ), .QN(n2971) );
  DFFARX1 \regfile_reg[9][2]  ( .D(n419), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[9][2] ), .QN(n3230) );
  DFFARX1 \regfile_reg[10][2]  ( .D(n418), .CLK(clk), .RSTB(n3758), .Q(
        \regfile[10][2] ), .QN(n3218) );
  DFFASX1 \regfile_reg[11][2]  ( .D(n417), .CLK(clk), .SETB(n3765), .Q(
        \regfile[11][2] ), .QN(n3466) );
  DFFASX1 \regfile_reg[12][2]  ( .D(n416), .CLK(clk), .SETB(n3764), .Q(
        \regfile[12][2] ), .QN(n3091) );
  DFFASX1 \regfile_reg[13][2]  ( .D(n415), .CLK(clk), .SETB(n3765), .Q(
        \regfile[13][2] ), .QN(n3350) );
  DFFASX1 \regfile_reg[14][2]  ( .D(n414), .CLK(clk), .SETB(n3765), .Q(
        \regfile[14][2] ), .QN(n3478) );
  DFFARX1 \regfile_reg[15][2]  ( .D(n413), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[15][2] ), .QN(n3103) );
  DFFARX1 \regfile_reg[0][1]  ( .D(n412), .CLK(clk), .RSTB(n3756), .Q(
        \regfile[0][1] ), .QN(n2970) );
  DFFASX1 \regfile_reg[1][1]  ( .D(n411), .CLK(clk), .SETB(n3765), .Q(
        \regfile[1][1] ), .QN(n3349) );
  DFFASX1 \regfile_reg[2][1]  ( .D(n410), .CLK(clk), .SETB(n3765), .Q(
        \regfile[2][1] ), .QN(n3477) );
  DFFARX1 \regfile_reg[3][1]  ( .D(n409), .CLK(clk), .RSTB(n3745), .Q(
        \regfile[3][1] ), .QN(n3102) );
  DFFARX1 \regfile_reg[4][1]  ( .D(n408), .CLK(clk), .RSTB(n3743), .Q(
        \regfile[4][1] ), .QN(n2969) );
  DFFASX1 \regfile_reg[5][1]  ( .D(n407), .CLK(clk), .SETB(n3765), .Q(
        \regfile[5][1] ), .QN(n3348) );
  DFFASX1 \regfile_reg[6][1]  ( .D(n406), .CLK(clk), .SETB(n3764), .Q(
        \regfile[6][1] ), .QN(n3476) );
  DFFARX1 \regfile_reg[7][1]  ( .D(n405), .CLK(clk), .RSTB(n3739), .Q(
        \regfile[7][1] ), .QN(n3101) );
  DFFARX1 \regfile_reg[8][1]  ( .D(n404), .CLK(clk), .RSTB(n3738), .Q(
        \regfile[8][1] ), .QN(n2968) );
  DFFASX1 \regfile_reg[9][1]  ( .D(n403), .CLK(clk), .SETB(n3764), .Q(
        \regfile[9][1] ), .QN(n3347) );
  DFFASX1 \regfile_reg[10][1]  ( .D(n402), .CLK(clk), .SETB(n3764), .Q(
        \regfile[10][1] ), .QN(n3475) );
  DFFARX1 \regfile_reg[11][1]  ( .D(n401), .CLK(clk), .RSTB(n3733), .Q(
        \regfile[11][1] ), .QN(n3100) );
  DFFARX1 \regfile_reg[12][1]  ( .D(n400), .CLK(clk), .RSTB(n3749), .Q(
        \regfile[12][1] ), .QN(n2967) );
  DFFASX1 \regfile_reg[13][1]  ( .D(n399), .CLK(clk), .SETB(n3764), .Q(
        \regfile[13][1] ), .QN(n3346) );
  DFFASX1 \regfile_reg[14][1]  ( .D(n398), .CLK(clk), .SETB(n3764), .Q(
        \regfile[14][1] ), .QN(n3474) );
  DFFARX1 \regfile_reg[15][1]  ( .D(n397), .CLK(clk), .RSTB(n3751), .Q(
        \regfile[15][1] ), .QN(n3099) );
  DFFASX1 \regfile_reg[0][0]  ( .D(n396), .CLK(clk), .SETB(n3764), .Q(
        \regfile[0][0] ), .QN(n3090) );
  DFFARX1 \regfile_reg[1][0]  ( .D(n395), .CLK(clk), .RSTB(n3746), .Q(
        \regfile[1][0] ), .QN(n3229) );
  DFFASX1 \regfile_reg[2][0]  ( .D(n394), .CLK(clk), .SETB(n3764), .Q(
        \regfile[2][0] ), .QN(n3473) );
  DFFARX1 \regfile_reg[3][0]  ( .D(n393), .CLK(clk), .RSTB(n3724), .Q(
        \regfile[3][0] ), .QN(n3098) );
  DFFASX1 \regfile_reg[4][0]  ( .D(n392), .CLK(clk), .SETB(n3763), .Q(
        \regfile[4][0] ), .QN(n3089) );
  DFFARX1 \regfile_reg[5][0]  ( .D(n391), .CLK(clk), .RSTB(n3727), .Q(
        \regfile[5][0] ), .QN(n3228) );
  DFFASX1 \regfile_reg[6][0]  ( .D(n390), .CLK(clk), .SETB(n3764), .Q(
        \regfile[6][0] ), .QN(n3472) );
  DFFARX1 \regfile_reg[7][0]  ( .D(n389), .CLK(clk), .RSTB(n3729), .Q(
        \regfile[7][0] ), .QN(n3097) );
  DFFASX1 \regfile_reg[8][0]  ( .D(n388), .CLK(clk), .SETB(n3763), .Q(
        \regfile[8][0] ), .QN(n3088) );
  DFFARX1 \regfile_reg[9][0]  ( .D(n387), .CLK(clk), .RSTB(n3732), .Q(
        \regfile[9][0] ), .QN(n3227) );
  DFFASX1 \regfile_reg[10][0]  ( .D(n386), .CLK(clk), .SETB(n3765), .Q(
        \regfile[10][0] ), .QN(n3471) );
  DFFARX1 \regfile_reg[11][0]  ( .D(n385), .CLK(clk), .RSTB(n3759), .Q(
        \regfile[11][0] ), .QN(n3096) );
  DFFASX1 \regfile_reg[12][0]  ( .D(n384), .CLK(clk), .SETB(n3765), .Q(
        \regfile[12][0] ), .QN(n3087) );
  DFFARX1 \regfile_reg[13][0]  ( .D(n383), .CLK(clk), .RSTB(n3761), .Q(
        \regfile[13][0] ), .QN(n3226) );
  DFFASX1 \regfile_reg[14][0]  ( .D(n382), .CLK(clk), .SETB(n3765), .Q(
        \regfile[14][0] ), .QN(n3470) );
  DFFARX1 \regfile_reg[15][0]  ( .D(n381), .CLK(clk), .RSTB(n3755), .Q(
        \regfile[15][0] ), .QN(n3095) );
  AO22X1 U1644 ( .IN1(n3810), .IN2(n3772), .IN3(n3768), .IN4(n2199), .Q(n964)
         );
  NAND4X0 U1645 ( .IN1(n2200), .IN2(n2201), .IN3(n2202), .IN4(n2203), .QN(
        n2199) );
  OA221X1 U1646 ( .IN1(n3721), .IN2(n3217), .IN3(n3718), .IN4(n3465), .IN5(
        n2206), .Q(n2203) );
  OA22X1 U1647 ( .IN1(n3715), .IN2(n3086), .IN3(n3712), .IN4(n3345), .Q(n2206)
         );
  OA221X1 U1648 ( .IN1(n3709), .IN2(n3216), .IN3(n3706), .IN4(n3464), .IN5(
        n2211), .Q(n2202) );
  OA22X1 U1649 ( .IN1(n3703), .IN2(n3085), .IN3(n3700), .IN4(n3344), .Q(n2211)
         );
  OA221X1 U1650 ( .IN1(n3697), .IN2(n3215), .IN3(n3694), .IN4(n3463), .IN5(
        n2216), .Q(n2201) );
  OA22X1 U1651 ( .IN1(n3691), .IN2(n3084), .IN3(n3688), .IN4(n3343), .Q(n2216)
         );
  OA221X1 U1652 ( .IN1(n3685), .IN2(n3214), .IN3(n3682), .IN4(n3462), .IN5(
        n2221), .Q(n2200) );
  OA22X1 U1653 ( .IN1(n3679), .IN2(n3083), .IN3(n3676), .IN4(n3342), .Q(n2221)
         );
  AO22X1 U1654 ( .IN1(IFID_B[30]), .IN2(n3772), .IN3(n3768), .IN4(n2224), .Q(
        n963) );
  NAND4X0 U1655 ( .IN1(n2225), .IN2(n2226), .IN3(n2227), .IN4(n2228), .QN(
        n2224) );
  OA221X1 U1656 ( .IN1(n3721), .IN2(n3213), .IN3(n3718), .IN4(n3461), .IN5(
        n2229), .Q(n2228) );
  OA22X1 U1657 ( .IN1(n3715), .IN2(n3082), .IN3(n3712), .IN4(n3341), .Q(n2229)
         );
  OA221X1 U1658 ( .IN1(n3709), .IN2(n3212), .IN3(n3706), .IN4(n3460), .IN5(
        n2230), .Q(n2227) );
  OA22X1 U1659 ( .IN1(n3703), .IN2(n3081), .IN3(n3700), .IN4(n3340), .Q(n2230)
         );
  OA221X1 U1660 ( .IN1(n3697), .IN2(n3211), .IN3(n3694), .IN4(n3459), .IN5(
        n2231), .Q(n2226) );
  OA22X1 U1661 ( .IN1(n3691), .IN2(n3080), .IN3(n3688), .IN4(n3339), .Q(n2231)
         );
  OA221X1 U1662 ( .IN1(n3685), .IN2(n3210), .IN3(n3682), .IN4(n3458), .IN5(
        n2232), .Q(n2225) );
  OA22X1 U1663 ( .IN1(n3679), .IN2(n3079), .IN3(n3676), .IN4(n3338), .Q(n2232)
         );
  AO22X1 U1664 ( .IN1(IFID_B[29]), .IN2(n3772), .IN3(n3768), .IN4(n2233), .Q(
        n962) );
  NAND4X0 U1665 ( .IN1(n2234), .IN2(n2235), .IN3(n2236), .IN4(n2237), .QN(
        n2233) );
  OA221X1 U1666 ( .IN1(n3721), .IN2(n3209), .IN3(n3718), .IN4(n3457), .IN5(
        n2238), .Q(n2237) );
  OA22X1 U1667 ( .IN1(n3715), .IN2(n3078), .IN3(n3712), .IN4(n3337), .Q(n2238)
         );
  OA221X1 U1668 ( .IN1(n3709), .IN2(n3208), .IN3(n3706), .IN4(n3456), .IN5(
        n2239), .Q(n2236) );
  OA22X1 U1669 ( .IN1(n3703), .IN2(n3077), .IN3(n3700), .IN4(n3336), .Q(n2239)
         );
  OA221X1 U1670 ( .IN1(n3697), .IN2(n3207), .IN3(n3694), .IN4(n3455), .IN5(
        n2240), .Q(n2235) );
  OA22X1 U1671 ( .IN1(n3691), .IN2(n3076), .IN3(n3688), .IN4(n3335), .Q(n2240)
         );
  OA221X1 U1672 ( .IN1(n3685), .IN2(n3206), .IN3(n3682), .IN4(n3454), .IN5(
        n2241), .Q(n2234) );
  OA22X1 U1673 ( .IN1(n3679), .IN2(n3075), .IN3(n3676), .IN4(n3334), .Q(n2241)
         );
  AO22X1 U1674 ( .IN1(IFID_B[28]), .IN2(n3772), .IN3(n3768), .IN4(n2242), .Q(
        n961) );
  NAND4X0 U1675 ( .IN1(n2243), .IN2(n2244), .IN3(n2245), .IN4(n2246), .QN(
        n2242) );
  OA221X1 U1676 ( .IN1(n3721), .IN2(n3205), .IN3(n3718), .IN4(n3453), .IN5(
        n2247), .Q(n2246) );
  OA22X1 U1677 ( .IN1(n3715), .IN2(n3074), .IN3(n3712), .IN4(n3333), .Q(n2247)
         );
  OA221X1 U1678 ( .IN1(n3709), .IN2(n3204), .IN3(n3706), .IN4(n3452), .IN5(
        n2248), .Q(n2245) );
  OA22X1 U1679 ( .IN1(n3703), .IN2(n3073), .IN3(n3700), .IN4(n3332), .Q(n2248)
         );
  OA221X1 U1680 ( .IN1(n3697), .IN2(n3203), .IN3(n3694), .IN4(n3451), .IN5(
        n2249), .Q(n2244) );
  OA22X1 U1681 ( .IN1(n3691), .IN2(n3072), .IN3(n3688), .IN4(n3331), .Q(n2249)
         );
  OA221X1 U1682 ( .IN1(n3685), .IN2(n3202), .IN3(n3682), .IN4(n3450), .IN5(
        n2250), .Q(n2243) );
  OA22X1 U1683 ( .IN1(n3679), .IN2(n3071), .IN3(n3676), .IN4(n3330), .Q(n2250)
         );
  AO22X1 U1684 ( .IN1(IFID_B[27]), .IN2(n3773), .IN3(n3768), .IN4(n2251), .Q(
        n960) );
  NAND4X0 U1685 ( .IN1(n2252), .IN2(n2253), .IN3(n2254), .IN4(n2255), .QN(
        n2251) );
  OA221X1 U1686 ( .IN1(n3721), .IN2(n3201), .IN3(n3718), .IN4(n3449), .IN5(
        n2256), .Q(n2255) );
  OA22X1 U1687 ( .IN1(n3715), .IN2(n3070), .IN3(n3712), .IN4(n3329), .Q(n2256)
         );
  OA221X1 U1688 ( .IN1(n3709), .IN2(n3200), .IN3(n3706), .IN4(n3448), .IN5(
        n2257), .Q(n2254) );
  OA22X1 U1689 ( .IN1(n3703), .IN2(n3069), .IN3(n3700), .IN4(n3328), .Q(n2257)
         );
  OA221X1 U1690 ( .IN1(n3697), .IN2(n3199), .IN3(n3694), .IN4(n3447), .IN5(
        n2258), .Q(n2253) );
  OA22X1 U1691 ( .IN1(n3691), .IN2(n3068), .IN3(n3688), .IN4(n3327), .Q(n2258)
         );
  OA221X1 U1692 ( .IN1(n3685), .IN2(n3198), .IN3(n3682), .IN4(n3446), .IN5(
        n2259), .Q(n2252) );
  OA22X1 U1693 ( .IN1(n3679), .IN2(n3067), .IN3(n3676), .IN4(n3326), .Q(n2259)
         );
  AO22X1 U1694 ( .IN1(IFID_B[26]), .IN2(n3773), .IN3(n3768), .IN4(n2260), .Q(
        n959) );
  NAND4X0 U1695 ( .IN1(n2261), .IN2(n2262), .IN3(n2263), .IN4(n2264), .QN(
        n2260) );
  OA221X1 U1696 ( .IN1(n3721), .IN2(n3197), .IN3(n3718), .IN4(n3445), .IN5(
        n2265), .Q(n2264) );
  OA22X1 U1697 ( .IN1(n3715), .IN2(n3066), .IN3(n3712), .IN4(n3325), .Q(n2265)
         );
  OA221X1 U1698 ( .IN1(n3709), .IN2(n3196), .IN3(n3706), .IN4(n3444), .IN5(
        n2266), .Q(n2263) );
  OA22X1 U1699 ( .IN1(n3703), .IN2(n3065), .IN3(n3700), .IN4(n3324), .Q(n2266)
         );
  OA221X1 U1700 ( .IN1(n3697), .IN2(n3195), .IN3(n3694), .IN4(n3443), .IN5(
        n2267), .Q(n2262) );
  OA22X1 U1701 ( .IN1(n3691), .IN2(n3064), .IN3(n3688), .IN4(n3323), .Q(n2267)
         );
  OA221X1 U1702 ( .IN1(n3685), .IN2(n3194), .IN3(n3682), .IN4(n3442), .IN5(
        n2268), .Q(n2261) );
  OA22X1 U1703 ( .IN1(n3679), .IN2(n3063), .IN3(n3676), .IN4(n3322), .Q(n2268)
         );
  AO22X1 U1704 ( .IN1(IFID_B[25]), .IN2(n3773), .IN3(n3768), .IN4(n2269), .Q(
        n958) );
  NAND4X0 U1705 ( .IN1(n2270), .IN2(n2271), .IN3(n2272), .IN4(n2273), .QN(
        n2269) );
  OA221X1 U1706 ( .IN1(n3721), .IN2(n3193), .IN3(n3718), .IN4(n3441), .IN5(
        n2274), .Q(n2273) );
  OA22X1 U1707 ( .IN1(n3715), .IN2(n3062), .IN3(n3712), .IN4(n3321), .Q(n2274)
         );
  OA221X1 U1708 ( .IN1(n3709), .IN2(n3192), .IN3(n3706), .IN4(n3440), .IN5(
        n2275), .Q(n2272) );
  OA22X1 U1709 ( .IN1(n3703), .IN2(n3061), .IN3(n3700), .IN4(n3320), .Q(n2275)
         );
  OA221X1 U1710 ( .IN1(n3697), .IN2(n3191), .IN3(n3694), .IN4(n3439), .IN5(
        n2276), .Q(n2271) );
  OA22X1 U1711 ( .IN1(n3691), .IN2(n3060), .IN3(n3688), .IN4(n3319), .Q(n2276)
         );
  OA221X1 U1712 ( .IN1(n3685), .IN2(n3190), .IN3(n3682), .IN4(n3438), .IN5(
        n2277), .Q(n2270) );
  OA22X1 U1713 ( .IN1(n3679), .IN2(n3059), .IN3(n3676), .IN4(n3318), .Q(n2277)
         );
  AO22X1 U1714 ( .IN1(IFID_B[24]), .IN2(n3773), .IN3(n3768), .IN4(n2278), .Q(
        n957) );
  NAND4X0 U1715 ( .IN1(n2279), .IN2(n2280), .IN3(n2281), .IN4(n2282), .QN(
        n2278) );
  OA221X1 U1716 ( .IN1(n3721), .IN2(n3189), .IN3(n3718), .IN4(n3437), .IN5(
        n2283), .Q(n2282) );
  OA22X1 U1717 ( .IN1(n3715), .IN2(n3058), .IN3(n3712), .IN4(n3317), .Q(n2283)
         );
  OA221X1 U1718 ( .IN1(n3709), .IN2(n3188), .IN3(n3706), .IN4(n3436), .IN5(
        n2284), .Q(n2281) );
  OA22X1 U1719 ( .IN1(n3703), .IN2(n3057), .IN3(n3700), .IN4(n3316), .Q(n2284)
         );
  OA221X1 U1720 ( .IN1(n3697), .IN2(n3187), .IN3(n3694), .IN4(n3435), .IN5(
        n2285), .Q(n2280) );
  OA22X1 U1721 ( .IN1(n3691), .IN2(n3056), .IN3(n3688), .IN4(n3315), .Q(n2285)
         );
  OA221X1 U1722 ( .IN1(n3685), .IN2(n3186), .IN3(n3682), .IN4(n3434), .IN5(
        n2286), .Q(n2279) );
  OA22X1 U1723 ( .IN1(n3679), .IN2(n3055), .IN3(n3676), .IN4(n3314), .Q(n2286)
         );
  AO22X1 U1724 ( .IN1(IFID_B[23]), .IN2(n3773), .IN3(n3768), .IN4(n2287), .Q(
        n956) );
  NAND4X0 U1725 ( .IN1(n2288), .IN2(n2289), .IN3(n2290), .IN4(n2291), .QN(
        n2287) );
  OA221X1 U1726 ( .IN1(n3721), .IN2(n3185), .IN3(n3718), .IN4(n3433), .IN5(
        n2292), .Q(n2291) );
  OA22X1 U1727 ( .IN1(n3715), .IN2(n3054), .IN3(n3712), .IN4(n3313), .Q(n2292)
         );
  OA221X1 U1728 ( .IN1(n3709), .IN2(n3184), .IN3(n3706), .IN4(n3432), .IN5(
        n2293), .Q(n2290) );
  OA22X1 U1729 ( .IN1(n3703), .IN2(n3053), .IN3(n3700), .IN4(n3312), .Q(n2293)
         );
  OA221X1 U1730 ( .IN1(n3697), .IN2(n3183), .IN3(n3694), .IN4(n3431), .IN5(
        n2294), .Q(n2289) );
  OA22X1 U1731 ( .IN1(n3691), .IN2(n3052), .IN3(n3688), .IN4(n3311), .Q(n2294)
         );
  OA221X1 U1732 ( .IN1(n3685), .IN2(n3182), .IN3(n3682), .IN4(n3430), .IN5(
        n2295), .Q(n2288) );
  OA22X1 U1733 ( .IN1(n3679), .IN2(n3051), .IN3(n3676), .IN4(n3310), .Q(n2295)
         );
  AO22X1 U1734 ( .IN1(IFID_B[22]), .IN2(n3773), .IN3(n3768), .IN4(n2296), .Q(
        n955) );
  NAND4X0 U1735 ( .IN1(n2297), .IN2(n2298), .IN3(n2299), .IN4(n2300), .QN(
        n2296) );
  OA221X1 U1736 ( .IN1(n3721), .IN2(n3181), .IN3(n3718), .IN4(n3429), .IN5(
        n2301), .Q(n2300) );
  OA22X1 U1737 ( .IN1(n3715), .IN2(n3050), .IN3(n3712), .IN4(n3309), .Q(n2301)
         );
  OA221X1 U1738 ( .IN1(n3709), .IN2(n3180), .IN3(n3706), .IN4(n3428), .IN5(
        n2302), .Q(n2299) );
  OA22X1 U1739 ( .IN1(n3703), .IN2(n3049), .IN3(n3700), .IN4(n3308), .Q(n2302)
         );
  OA221X1 U1740 ( .IN1(n3697), .IN2(n3179), .IN3(n3694), .IN4(n3427), .IN5(
        n2303), .Q(n2298) );
  OA22X1 U1741 ( .IN1(n3691), .IN2(n3048), .IN3(n3688), .IN4(n3307), .Q(n2303)
         );
  OA221X1 U1742 ( .IN1(n3685), .IN2(n3178), .IN3(n3682), .IN4(n3426), .IN5(
        n2304), .Q(n2297) );
  OA22X1 U1743 ( .IN1(n3679), .IN2(n3047), .IN3(n3676), .IN4(n3306), .Q(n2304)
         );
  AO22X1 U1744 ( .IN1(IFID_B[21]), .IN2(n3773), .IN3(n3768), .IN4(n2305), .Q(
        n954) );
  NAND4X0 U1745 ( .IN1(n2306), .IN2(n2307), .IN3(n2308), .IN4(n2309), .QN(
        n2305) );
  OA221X1 U1746 ( .IN1(n3721), .IN2(n3177), .IN3(n3718), .IN4(n3425), .IN5(
        n2310), .Q(n2309) );
  OA22X1 U1747 ( .IN1(n3715), .IN2(n3046), .IN3(n3712), .IN4(n3305), .Q(n2310)
         );
  OA221X1 U1748 ( .IN1(n3709), .IN2(n3176), .IN3(n3706), .IN4(n3424), .IN5(
        n2311), .Q(n2308) );
  OA22X1 U1749 ( .IN1(n3703), .IN2(n3045), .IN3(n3700), .IN4(n3304), .Q(n2311)
         );
  OA221X1 U1750 ( .IN1(n3697), .IN2(n3175), .IN3(n3694), .IN4(n3423), .IN5(
        n2312), .Q(n2307) );
  OA22X1 U1751 ( .IN1(n3691), .IN2(n3044), .IN3(n3688), .IN4(n3303), .Q(n2312)
         );
  OA221X1 U1752 ( .IN1(n3685), .IN2(n3174), .IN3(n3682), .IN4(n3422), .IN5(
        n2313), .Q(n2306) );
  OA22X1 U1753 ( .IN1(n3679), .IN2(n3043), .IN3(n3676), .IN4(n3302), .Q(n2313)
         );
  AO22X1 U1754 ( .IN1(IFID_B[20]), .IN2(n3773), .IN3(n3767), .IN4(n2314), .Q(
        n953) );
  NAND4X0 U1755 ( .IN1(n2315), .IN2(n2316), .IN3(n2317), .IN4(n2318), .QN(
        n2314) );
  OA221X1 U1756 ( .IN1(n3721), .IN2(n3173), .IN3(n3718), .IN4(n3421), .IN5(
        n2319), .Q(n2318) );
  OA22X1 U1757 ( .IN1(n3715), .IN2(n3042), .IN3(n3712), .IN4(n3301), .Q(n2319)
         );
  OA221X1 U1758 ( .IN1(n3709), .IN2(n3172), .IN3(n3706), .IN4(n3420), .IN5(
        n2320), .Q(n2317) );
  OA22X1 U1759 ( .IN1(n3703), .IN2(n3041), .IN3(n3700), .IN4(n3300), .Q(n2320)
         );
  OA221X1 U1760 ( .IN1(n3697), .IN2(n3171), .IN3(n3694), .IN4(n3419), .IN5(
        n2321), .Q(n2316) );
  OA22X1 U1761 ( .IN1(n3691), .IN2(n3040), .IN3(n3688), .IN4(n3299), .Q(n2321)
         );
  OA221X1 U1762 ( .IN1(n3685), .IN2(n3170), .IN3(n3682), .IN4(n3418), .IN5(
        n2322), .Q(n2315) );
  OA22X1 U1763 ( .IN1(n3679), .IN2(n3039), .IN3(n3676), .IN4(n3298), .Q(n2322)
         );
  AO22X1 U1764 ( .IN1(IFID_B[19]), .IN2(n3773), .IN3(n3767), .IN4(n2323), .Q(
        n952) );
  NAND4X0 U1765 ( .IN1(n2324), .IN2(n2325), .IN3(n2326), .IN4(n2327), .QN(
        n2323) );
  OA221X1 U1766 ( .IN1(n3722), .IN2(n3169), .IN3(n3719), .IN4(n3417), .IN5(
        n2328), .Q(n2327) );
  OA22X1 U1767 ( .IN1(n3716), .IN2(n3038), .IN3(n3713), .IN4(n3297), .Q(n2328)
         );
  OA221X1 U1768 ( .IN1(n3710), .IN2(n3168), .IN3(n3707), .IN4(n3416), .IN5(
        n2329), .Q(n2326) );
  OA22X1 U1769 ( .IN1(n3704), .IN2(n3037), .IN3(n3701), .IN4(n3296), .Q(n2329)
         );
  OA221X1 U1770 ( .IN1(n3698), .IN2(n3167), .IN3(n3695), .IN4(n3415), .IN5(
        n2330), .Q(n2325) );
  OA22X1 U1771 ( .IN1(n3692), .IN2(n3036), .IN3(n3689), .IN4(n3295), .Q(n2330)
         );
  OA221X1 U1772 ( .IN1(n3686), .IN2(n3166), .IN3(n3683), .IN4(n3414), .IN5(
        n2331), .Q(n2324) );
  OA22X1 U1773 ( .IN1(n3680), .IN2(n3035), .IN3(n3677), .IN4(n3294), .Q(n2331)
         );
  AO22X1 U1774 ( .IN1(IFID_B[18]), .IN2(n3773), .IN3(n3767), .IN4(n2332), .Q(
        n951) );
  NAND4X0 U1775 ( .IN1(n2333), .IN2(n2334), .IN3(n2335), .IN4(n2336), .QN(
        n2332) );
  OA221X1 U1776 ( .IN1(n3722), .IN2(n3165), .IN3(n3719), .IN4(n3413), .IN5(
        n2337), .Q(n2336) );
  OA22X1 U1777 ( .IN1(n3716), .IN2(n3034), .IN3(n3713), .IN4(n3293), .Q(n2337)
         );
  OA221X1 U1778 ( .IN1(n3710), .IN2(n3164), .IN3(n3707), .IN4(n3412), .IN5(
        n2338), .Q(n2335) );
  OA22X1 U1779 ( .IN1(n3704), .IN2(n3033), .IN3(n3701), .IN4(n3292), .Q(n2338)
         );
  OA221X1 U1780 ( .IN1(n3698), .IN2(n3163), .IN3(n3695), .IN4(n3411), .IN5(
        n2339), .Q(n2334) );
  OA22X1 U1781 ( .IN1(n3692), .IN2(n3032), .IN3(n3689), .IN4(n3291), .Q(n2339)
         );
  OA221X1 U1782 ( .IN1(n3686), .IN2(n3162), .IN3(n3683), .IN4(n3410), .IN5(
        n2340), .Q(n2333) );
  OA22X1 U1783 ( .IN1(n3680), .IN2(n3031), .IN3(n3677), .IN4(n3290), .Q(n2340)
         );
  AO22X1 U1784 ( .IN1(IFID_B[17]), .IN2(n3773), .IN3(n3767), .IN4(n2341), .Q(
        n950) );
  NAND4X0 U1785 ( .IN1(n2342), .IN2(n2343), .IN3(n2344), .IN4(n2345), .QN(
        n2341) );
  OA221X1 U1786 ( .IN1(n3722), .IN2(n3161), .IN3(n3719), .IN4(n3409), .IN5(
        n2346), .Q(n2345) );
  OA22X1 U1787 ( .IN1(n3716), .IN2(n3030), .IN3(n3713), .IN4(n3289), .Q(n2346)
         );
  OA221X1 U1788 ( .IN1(n3710), .IN2(n3160), .IN3(n3707), .IN4(n3408), .IN5(
        n2347), .Q(n2344) );
  OA22X1 U1789 ( .IN1(n3704), .IN2(n3029), .IN3(n3701), .IN4(n3288), .Q(n2347)
         );
  OA221X1 U1790 ( .IN1(n3698), .IN2(n3159), .IN3(n3695), .IN4(n3407), .IN5(
        n2348), .Q(n2343) );
  OA22X1 U1791 ( .IN1(n3692), .IN2(n3028), .IN3(n3689), .IN4(n3287), .Q(n2348)
         );
  OA221X1 U1792 ( .IN1(n3686), .IN2(n3158), .IN3(n3683), .IN4(n3406), .IN5(
        n2349), .Q(n2342) );
  OA22X1 U1793 ( .IN1(n3680), .IN2(n3027), .IN3(n3677), .IN4(n3286), .Q(n2349)
         );
  AO22X1 U1794 ( .IN1(IFID_B[16]), .IN2(n3773), .IN3(n3767), .IN4(n2350), .Q(
        n949) );
  NAND4X0 U1795 ( .IN1(n2351), .IN2(n2352), .IN3(n2353), .IN4(n2354), .QN(
        n2350) );
  OA221X1 U1796 ( .IN1(n3722), .IN2(n3157), .IN3(n3719), .IN4(n3405), .IN5(
        n2355), .Q(n2354) );
  OA22X1 U1797 ( .IN1(n3716), .IN2(n3026), .IN3(n3713), .IN4(n3285), .Q(n2355)
         );
  OA221X1 U1798 ( .IN1(n3710), .IN2(n3156), .IN3(n3707), .IN4(n3404), .IN5(
        n2356), .Q(n2353) );
  OA22X1 U1799 ( .IN1(n3704), .IN2(n3025), .IN3(n3701), .IN4(n3284), .Q(n2356)
         );
  OA221X1 U1800 ( .IN1(n3698), .IN2(n3155), .IN3(n3695), .IN4(n3403), .IN5(
        n2357), .Q(n2352) );
  OA22X1 U1801 ( .IN1(n3692), .IN2(n3024), .IN3(n3689), .IN4(n3283), .Q(n2357)
         );
  OA221X1 U1802 ( .IN1(n3686), .IN2(n3154), .IN3(n3683), .IN4(n3402), .IN5(
        n2358), .Q(n2351) );
  OA22X1 U1803 ( .IN1(n3680), .IN2(n3023), .IN3(n3677), .IN4(n3282), .Q(n2358)
         );
  AO22X1 U1804 ( .IN1(IFID_B[15]), .IN2(n3773), .IN3(n3767), .IN4(n2359), .Q(
        n948) );
  NAND4X0 U1805 ( .IN1(n2360), .IN2(n2361), .IN3(n2362), .IN4(n2363), .QN(
        n2359) );
  OA221X1 U1806 ( .IN1(n3722), .IN2(n3153), .IN3(n3719), .IN4(n3401), .IN5(
        n2364), .Q(n2363) );
  OA22X1 U1807 ( .IN1(n3716), .IN2(n3022), .IN3(n3713), .IN4(n3281), .Q(n2364)
         );
  OA221X1 U1808 ( .IN1(n3710), .IN2(n3152), .IN3(n3707), .IN4(n3400), .IN5(
        n2365), .Q(n2362) );
  OA22X1 U1809 ( .IN1(n3704), .IN2(n3021), .IN3(n3701), .IN4(n3280), .Q(n2365)
         );
  OA221X1 U1810 ( .IN1(n3698), .IN2(n3151), .IN3(n3695), .IN4(n3399), .IN5(
        n2366), .Q(n2361) );
  OA22X1 U1811 ( .IN1(n3692), .IN2(n3020), .IN3(n3689), .IN4(n3279), .Q(n2366)
         );
  OA221X1 U1812 ( .IN1(n3686), .IN2(n3150), .IN3(n3683), .IN4(n3398), .IN5(
        n2367), .Q(n2360) );
  OA22X1 U1813 ( .IN1(n3680), .IN2(n3019), .IN3(n3677), .IN4(n3278), .Q(n2367)
         );
  AO22X1 U1814 ( .IN1(IFID_B[14]), .IN2(n3773), .IN3(n3767), .IN4(n2368), .Q(
        n947) );
  NAND4X0 U1815 ( .IN1(n2369), .IN2(n2370), .IN3(n2371), .IN4(n2372), .QN(
        n2368) );
  OA221X1 U1816 ( .IN1(n3722), .IN2(n3149), .IN3(n3719), .IN4(n3397), .IN5(
        n2373), .Q(n2372) );
  OA22X1 U1817 ( .IN1(n3716), .IN2(n3018), .IN3(n3713), .IN4(n3277), .Q(n2373)
         );
  OA221X1 U1818 ( .IN1(n3710), .IN2(n3148), .IN3(n3707), .IN4(n3396), .IN5(
        n2374), .Q(n2371) );
  OA22X1 U1819 ( .IN1(n3704), .IN2(n3017), .IN3(n3701), .IN4(n3276), .Q(n2374)
         );
  OA221X1 U1820 ( .IN1(n3698), .IN2(n3147), .IN3(n3695), .IN4(n3395), .IN5(
        n2375), .Q(n2370) );
  OA22X1 U1821 ( .IN1(n3692), .IN2(n3016), .IN3(n3689), .IN4(n3275), .Q(n2375)
         );
  OA221X1 U1822 ( .IN1(n3686), .IN2(n3146), .IN3(n3683), .IN4(n3394), .IN5(
        n2376), .Q(n2369) );
  OA22X1 U1823 ( .IN1(n3680), .IN2(n3015), .IN3(n3677), .IN4(n3274), .Q(n2376)
         );
  AO22X1 U1824 ( .IN1(IFID_B[13]), .IN2(n3774), .IN3(n3767), .IN4(n2377), .Q(
        n946) );
  NAND4X0 U1825 ( .IN1(n2378), .IN2(n2379), .IN3(n2380), .IN4(n2381), .QN(
        n2377) );
  OA221X1 U1826 ( .IN1(n3722), .IN2(n3145), .IN3(n3719), .IN4(n3393), .IN5(
        n2382), .Q(n2381) );
  OA22X1 U1827 ( .IN1(n3716), .IN2(n3014), .IN3(n3713), .IN4(n3273), .Q(n2382)
         );
  OA221X1 U1828 ( .IN1(n3710), .IN2(n3144), .IN3(n3707), .IN4(n3392), .IN5(
        n2383), .Q(n2380) );
  OA22X1 U1829 ( .IN1(n3704), .IN2(n3013), .IN3(n3701), .IN4(n3272), .Q(n2383)
         );
  OA221X1 U1830 ( .IN1(n3698), .IN2(n3143), .IN3(n3695), .IN4(n3391), .IN5(
        n2384), .Q(n2379) );
  OA22X1 U1831 ( .IN1(n3692), .IN2(n3012), .IN3(n3689), .IN4(n3271), .Q(n2384)
         );
  OA221X1 U1832 ( .IN1(n3686), .IN2(n3142), .IN3(n3683), .IN4(n3390), .IN5(
        n2385), .Q(n2378) );
  OA22X1 U1833 ( .IN1(n3680), .IN2(n3011), .IN3(n3677), .IN4(n3270), .Q(n2385)
         );
  AO22X1 U1834 ( .IN1(IFID_B[12]), .IN2(n3774), .IN3(n3767), .IN4(n2386), .Q(
        n945) );
  NAND4X0 U1835 ( .IN1(n2387), .IN2(n2388), .IN3(n2389), .IN4(n2390), .QN(
        n2386) );
  OA221X1 U1836 ( .IN1(n3722), .IN2(n3141), .IN3(n3719), .IN4(n3389), .IN5(
        n2391), .Q(n2390) );
  OA22X1 U1837 ( .IN1(n3716), .IN2(n3010), .IN3(n3713), .IN4(n3269), .Q(n2391)
         );
  OA221X1 U1838 ( .IN1(n3710), .IN2(n3140), .IN3(n3707), .IN4(n3388), .IN5(
        n2392), .Q(n2389) );
  OA22X1 U1839 ( .IN1(n3704), .IN2(n3009), .IN3(n3701), .IN4(n3268), .Q(n2392)
         );
  OA221X1 U1840 ( .IN1(n3698), .IN2(n3139), .IN3(n3695), .IN4(n3387), .IN5(
        n2393), .Q(n2388) );
  OA22X1 U1841 ( .IN1(n3692), .IN2(n3008), .IN3(n3689), .IN4(n3267), .Q(n2393)
         );
  OA221X1 U1842 ( .IN1(n3686), .IN2(n3138), .IN3(n3683), .IN4(n3386), .IN5(
        n2394), .Q(n2387) );
  OA22X1 U1843 ( .IN1(n3680), .IN2(n3007), .IN3(n3677), .IN4(n3266), .Q(n2394)
         );
  AO22X1 U1844 ( .IN1(IFID_B[11]), .IN2(n3774), .IN3(n3767), .IN4(n2395), .Q(
        n944) );
  NAND4X0 U1845 ( .IN1(n2396), .IN2(n2397), .IN3(n2398), .IN4(n2399), .QN(
        n2395) );
  OA221X1 U1846 ( .IN1(n3722), .IN2(n3137), .IN3(n3719), .IN4(n3385), .IN5(
        n2400), .Q(n2399) );
  OA22X1 U1847 ( .IN1(n3716), .IN2(n3006), .IN3(n3713), .IN4(n3265), .Q(n2400)
         );
  OA221X1 U1848 ( .IN1(n3710), .IN2(n3136), .IN3(n3707), .IN4(n3384), .IN5(
        n2401), .Q(n2398) );
  OA22X1 U1849 ( .IN1(n3704), .IN2(n3005), .IN3(n3701), .IN4(n3264), .Q(n2401)
         );
  OA221X1 U1850 ( .IN1(n3698), .IN2(n3135), .IN3(n3695), .IN4(n3383), .IN5(
        n2402), .Q(n2397) );
  OA22X1 U1851 ( .IN1(n3692), .IN2(n3004), .IN3(n3689), .IN4(n3263), .Q(n2402)
         );
  OA221X1 U1852 ( .IN1(n3686), .IN2(n3134), .IN3(n3683), .IN4(n3382), .IN5(
        n2403), .Q(n2396) );
  OA22X1 U1853 ( .IN1(n3680), .IN2(n3003), .IN3(n3677), .IN4(n3262), .Q(n2403)
         );
  AO22X1 U1854 ( .IN1(IFID_B[10]), .IN2(n3774), .IN3(n3767), .IN4(n2404), .Q(
        n943) );
  NAND4X0 U1855 ( .IN1(n2405), .IN2(n2406), .IN3(n2407), .IN4(n2408), .QN(
        n2404) );
  OA221X1 U1856 ( .IN1(n3722), .IN2(n3133), .IN3(n3719), .IN4(n3381), .IN5(
        n2409), .Q(n2408) );
  OA22X1 U1857 ( .IN1(n3716), .IN2(n3002), .IN3(n3713), .IN4(n3261), .Q(n2409)
         );
  OA221X1 U1858 ( .IN1(n3710), .IN2(n3132), .IN3(n3707), .IN4(n3380), .IN5(
        n2410), .Q(n2407) );
  OA22X1 U1859 ( .IN1(n3704), .IN2(n3001), .IN3(n3701), .IN4(n3260), .Q(n2410)
         );
  OA221X1 U1860 ( .IN1(n3698), .IN2(n3131), .IN3(n3695), .IN4(n3379), .IN5(
        n2411), .Q(n2406) );
  OA22X1 U1861 ( .IN1(n3692), .IN2(n3000), .IN3(n3689), .IN4(n3259), .Q(n2411)
         );
  OA221X1 U1862 ( .IN1(n3686), .IN2(n3130), .IN3(n3683), .IN4(n3378), .IN5(
        n2412), .Q(n2405) );
  OA22X1 U1863 ( .IN1(n3680), .IN2(n2999), .IN3(n3677), .IN4(n3258), .Q(n2412)
         );
  AO22X1 U1864 ( .IN1(IFID_B[9]), .IN2(n3774), .IN3(n3767), .IN4(n2413), .Q(
        n942) );
  NAND4X0 U1865 ( .IN1(n2414), .IN2(n2415), .IN3(n2416), .IN4(n2417), .QN(
        n2413) );
  OA221X1 U1866 ( .IN1(n3722), .IN2(n3129), .IN3(n3719), .IN4(n3377), .IN5(
        n2418), .Q(n2417) );
  OA22X1 U1867 ( .IN1(n3716), .IN2(n2998), .IN3(n3713), .IN4(n3257), .Q(n2418)
         );
  OA221X1 U1868 ( .IN1(n3710), .IN2(n3128), .IN3(n3707), .IN4(n3376), .IN5(
        n2419), .Q(n2416) );
  OA22X1 U1869 ( .IN1(n3704), .IN2(n2997), .IN3(n3701), .IN4(n3256), .Q(n2419)
         );
  OA221X1 U1870 ( .IN1(n3698), .IN2(n3127), .IN3(n3695), .IN4(n3375), .IN5(
        n2420), .Q(n2415) );
  OA22X1 U1871 ( .IN1(n3692), .IN2(n2996), .IN3(n3689), .IN4(n3255), .Q(n2420)
         );
  OA221X1 U1872 ( .IN1(n3686), .IN2(n3126), .IN3(n3683), .IN4(n3374), .IN5(
        n2421), .Q(n2414) );
  OA22X1 U1873 ( .IN1(n3680), .IN2(n2995), .IN3(n3677), .IN4(n3254), .Q(n2421)
         );
  AO22X1 U1874 ( .IN1(IFID_B[8]), .IN2(n3774), .IN3(n3767), .IN4(n2422), .Q(
        n941) );
  NAND4X0 U1875 ( .IN1(n2423), .IN2(n2424), .IN3(n2425), .IN4(n2426), .QN(
        n2422) );
  OA221X1 U1876 ( .IN1(n3722), .IN2(n3125), .IN3(n3719), .IN4(n3373), .IN5(
        n2427), .Q(n2426) );
  OA22X1 U1877 ( .IN1(n3716), .IN2(n2994), .IN3(n3713), .IN4(n3253), .Q(n2427)
         );
  OA221X1 U1878 ( .IN1(n3710), .IN2(n3124), .IN3(n3707), .IN4(n3372), .IN5(
        n2428), .Q(n2425) );
  OA22X1 U1879 ( .IN1(n3704), .IN2(n2993), .IN3(n3701), .IN4(n3252), .Q(n2428)
         );
  OA221X1 U1880 ( .IN1(n3698), .IN2(n3123), .IN3(n3695), .IN4(n3371), .IN5(
        n2429), .Q(n2424) );
  OA22X1 U1881 ( .IN1(n3692), .IN2(n2992), .IN3(n3689), .IN4(n3251), .Q(n2429)
         );
  OA221X1 U1882 ( .IN1(n3686), .IN2(n3122), .IN3(n3683), .IN4(n3370), .IN5(
        n2430), .Q(n2423) );
  OA22X1 U1883 ( .IN1(n3680), .IN2(n2991), .IN3(n3677), .IN4(n3250), .Q(n2430)
         );
  AO22X1 U1884 ( .IN1(IFID_B[7]), .IN2(n3774), .IN3(n3767), .IN4(n2431), .Q(
        n940) );
  NAND4X0 U1885 ( .IN1(n2432), .IN2(n2433), .IN3(n2434), .IN4(n2435), .QN(
        n2431) );
  OA221X1 U1886 ( .IN1(n3723), .IN2(n3121), .IN3(n3720), .IN4(n3369), .IN5(
        n2436), .Q(n2435) );
  OA22X1 U1887 ( .IN1(n3717), .IN2(n2990), .IN3(n3714), .IN4(n3249), .Q(n2436)
         );
  OA221X1 U1888 ( .IN1(n3711), .IN2(n3120), .IN3(n3708), .IN4(n3368), .IN5(
        n2437), .Q(n2434) );
  OA22X1 U1889 ( .IN1(n3705), .IN2(n2989), .IN3(n3702), .IN4(n3248), .Q(n2437)
         );
  OA221X1 U1890 ( .IN1(n3699), .IN2(n3119), .IN3(n3696), .IN4(n3367), .IN5(
        n2438), .Q(n2433) );
  OA22X1 U1891 ( .IN1(n3693), .IN2(n2988), .IN3(n3690), .IN4(n3247), .Q(n2438)
         );
  OA221X1 U1892 ( .IN1(n3687), .IN2(n3118), .IN3(n3684), .IN4(n3366), .IN5(
        n2439), .Q(n2432) );
  OA22X1 U1893 ( .IN1(n3681), .IN2(n2987), .IN3(n3678), .IN4(n3246), .Q(n2439)
         );
  AO22X1 U1894 ( .IN1(IFID_B[6]), .IN2(n3774), .IN3(n3767), .IN4(n2440), .Q(
        n939) );
  NAND4X0 U1895 ( .IN1(n2441), .IN2(n2442), .IN3(n2443), .IN4(n2444), .QN(
        n2440) );
  OA221X1 U1896 ( .IN1(n3723), .IN2(n3117), .IN3(n3720), .IN4(n3365), .IN5(
        n2445), .Q(n2444) );
  OA22X1 U1897 ( .IN1(n3717), .IN2(n2986), .IN3(n3714), .IN4(n3245), .Q(n2445)
         );
  OA221X1 U1898 ( .IN1(n3711), .IN2(n3116), .IN3(n3708), .IN4(n3364), .IN5(
        n2446), .Q(n2443) );
  OA22X1 U1899 ( .IN1(n3705), .IN2(n2985), .IN3(n3702), .IN4(n3244), .Q(n2446)
         );
  OA221X1 U1900 ( .IN1(n3699), .IN2(n3115), .IN3(n3696), .IN4(n3363), .IN5(
        n2447), .Q(n2442) );
  OA22X1 U1901 ( .IN1(n3693), .IN2(n2984), .IN3(n3690), .IN4(n3243), .Q(n2447)
         );
  OA221X1 U1902 ( .IN1(n3687), .IN2(n3114), .IN3(n3684), .IN4(n3362), .IN5(
        n2448), .Q(n2441) );
  OA22X1 U1903 ( .IN1(n3681), .IN2(n2983), .IN3(n3678), .IN4(n3242), .Q(n2448)
         );
  AO22X1 U1904 ( .IN1(IFID_B[5]), .IN2(n3774), .IN3(n3767), .IN4(n2449), .Q(
        n938) );
  NAND4X0 U1905 ( .IN1(n2450), .IN2(n2451), .IN3(n2452), .IN4(n2453), .QN(
        n2449) );
  OA221X1 U1906 ( .IN1(n3723), .IN2(n3113), .IN3(n3720), .IN4(n3361), .IN5(
        n2454), .Q(n2453) );
  OA22X1 U1907 ( .IN1(n3717), .IN2(n2982), .IN3(n3714), .IN4(n3241), .Q(n2454)
         );
  OA221X1 U1908 ( .IN1(n3711), .IN2(n3112), .IN3(n3708), .IN4(n3360), .IN5(
        n2455), .Q(n2452) );
  OA22X1 U1909 ( .IN1(n3705), .IN2(n2981), .IN3(n3702), .IN4(n3240), .Q(n2455)
         );
  OA221X1 U1910 ( .IN1(n3699), .IN2(n3111), .IN3(n3696), .IN4(n3359), .IN5(
        n2456), .Q(n2451) );
  OA22X1 U1911 ( .IN1(n3693), .IN2(n2980), .IN3(n3690), .IN4(n3239), .Q(n2456)
         );
  OA221X1 U1912 ( .IN1(n3687), .IN2(n3110), .IN3(n3684), .IN4(n3358), .IN5(
        n2457), .Q(n2450) );
  OA22X1 U1913 ( .IN1(n3681), .IN2(n2979), .IN3(n3678), .IN4(n3238), .Q(n2457)
         );
  AO22X1 U1914 ( .IN1(IFID_B[4]), .IN2(n3774), .IN3(n3767), .IN4(n2458), .Q(
        n937) );
  NAND4X0 U1915 ( .IN1(n2459), .IN2(n2460), .IN3(n2461), .IN4(n2462), .QN(
        n2458) );
  OA221X1 U1916 ( .IN1(n3723), .IN2(n3109), .IN3(n3720), .IN4(n3357), .IN5(
        n2463), .Q(n2462) );
  OA22X1 U1917 ( .IN1(n3717), .IN2(n2978), .IN3(n3714), .IN4(n3237), .Q(n2463)
         );
  OA221X1 U1918 ( .IN1(n3711), .IN2(n3108), .IN3(n3708), .IN4(n3356), .IN5(
        n2464), .Q(n2461) );
  OA22X1 U1919 ( .IN1(n3705), .IN2(n2977), .IN3(n3702), .IN4(n3236), .Q(n2464)
         );
  OA221X1 U1920 ( .IN1(n3699), .IN2(n3107), .IN3(n3696), .IN4(n3355), .IN5(
        n2465), .Q(n2460) );
  OA22X1 U1921 ( .IN1(n3693), .IN2(n2976), .IN3(n3690), .IN4(n3235), .Q(n2465)
         );
  OA221X1 U1922 ( .IN1(n3687), .IN2(n3469), .IN3(n3684), .IN4(n3221), .IN5(
        n2466), .Q(n2459) );
  OA22X1 U1923 ( .IN1(n3681), .IN2(n2975), .IN3(n3678), .IN4(n3234), .Q(n2466)
         );
  AO22X1 U1924 ( .IN1(IFID_B[3]), .IN2(n3774), .IN3(n3767), .IN4(n2467), .Q(
        n936) );
  NAND4X0 U1925 ( .IN1(n2468), .IN2(n2469), .IN3(n2470), .IN4(n2471), .QN(
        n2467) );
  OA221X1 U1926 ( .IN1(n3723), .IN2(n3106), .IN3(n3720), .IN4(n3354), .IN5(
        n2472), .Q(n2471) );
  OA22X1 U1927 ( .IN1(n3717), .IN2(n2974), .IN3(n3714), .IN4(n3233), .Q(n2472)
         );
  OA221X1 U1928 ( .IN1(n3711), .IN2(n3468), .IN3(n3708), .IN4(n3220), .IN5(
        n2473), .Q(n2470) );
  OA22X1 U1929 ( .IN1(n3705), .IN2(n2973), .IN3(n3702), .IN4(n3232), .Q(n2473)
         );
  OA221X1 U1930 ( .IN1(n3699), .IN2(n3222), .IN3(n3696), .IN4(n3481), .IN5(
        n2474), .Q(n2469) );
  OA22X1 U1931 ( .IN1(n3693), .IN2(n3094), .IN3(n3690), .IN4(n3353), .Q(n2474)
         );
  OA221X1 U1932 ( .IN1(n3687), .IN2(n3105), .IN3(n3684), .IN4(n3480), .IN5(
        n2475), .Q(n2468) );
  OA22X1 U1933 ( .IN1(n3681), .IN2(n3093), .IN3(n3678), .IN4(n3352), .Q(n2475)
         );
  AO22X1 U1934 ( .IN1(IFID_B[2]), .IN2(n3774), .IN3(n3767), .IN4(n2476), .Q(
        n935) );
  NAND4X0 U1935 ( .IN1(n2477), .IN2(n2478), .IN3(n2479), .IN4(n2480), .QN(
        n2476) );
  OA221X1 U1936 ( .IN1(n3723), .IN2(n3467), .IN3(n3720), .IN4(n3219), .IN5(
        n2481), .Q(n2480) );
  OA22X1 U1937 ( .IN1(n3717), .IN2(n2972), .IN3(n3714), .IN4(n3231), .Q(n2481)
         );
  OA221X1 U1938 ( .IN1(n3711), .IN2(n3104), .IN3(n3708), .IN4(n3479), .IN5(
        n2482), .Q(n2479) );
  OA22X1 U1939 ( .IN1(n3705), .IN2(n3092), .IN3(n3702), .IN4(n3351), .Q(n2482)
         );
  OA221X1 U1940 ( .IN1(n3699), .IN2(n3466), .IN3(n3696), .IN4(n3218), .IN5(
        n2483), .Q(n2478) );
  OA22X1 U1941 ( .IN1(n3693), .IN2(n2971), .IN3(n3690), .IN4(n3230), .Q(n2483)
         );
  OA221X1 U1942 ( .IN1(n3687), .IN2(n3103), .IN3(n3684), .IN4(n3478), .IN5(
        n2484), .Q(n2477) );
  OA22X1 U1943 ( .IN1(n3681), .IN2(n3091), .IN3(n3678), .IN4(n3350), .Q(n2484)
         );
  AO22X1 U1944 ( .IN1(IFID_B[1]), .IN2(n3774), .IN3(n3767), .IN4(n2485), .Q(
        n934) );
  NAND4X0 U1945 ( .IN1(n2486), .IN2(n2487), .IN3(n2488), .IN4(n2489), .QN(
        n2485) );
  OA221X1 U1946 ( .IN1(n3723), .IN2(n3102), .IN3(n3720), .IN4(n3477), .IN5(
        n2490), .Q(n2489) );
  OA22X1 U1947 ( .IN1(n3717), .IN2(n2970), .IN3(n3714), .IN4(n3349), .Q(n2490)
         );
  OA221X1 U1948 ( .IN1(n3711), .IN2(n3101), .IN3(n3708), .IN4(n3476), .IN5(
        n2491), .Q(n2488) );
  OA22X1 U1949 ( .IN1(n3705), .IN2(n2969), .IN3(n3702), .IN4(n3348), .Q(n2491)
         );
  OA221X1 U1950 ( .IN1(n3699), .IN2(n3100), .IN3(n3696), .IN4(n3475), .IN5(
        n2492), .Q(n2487) );
  OA22X1 U1951 ( .IN1(n3693), .IN2(n2968), .IN3(n3690), .IN4(n3347), .Q(n2492)
         );
  OA221X1 U1952 ( .IN1(n3687), .IN2(n3099), .IN3(n3684), .IN4(n3474), .IN5(
        n2493), .Q(n2486) );
  OA22X1 U1953 ( .IN1(n3681), .IN2(n2967), .IN3(n3678), .IN4(n3346), .Q(n2493)
         );
  AO22X1 U1954 ( .IN1(IFID_B[0]), .IN2(n3774), .IN3(n3767), .IN4(n2494), .Q(
        n933) );
  NAND4X0 U1955 ( .IN1(n2495), .IN2(n2496), .IN3(n2497), .IN4(n2498), .QN(
        n2494) );
  OA221X1 U1956 ( .IN1(n3723), .IN2(n3098), .IN3(n3720), .IN4(n3473), .IN5(
        n2499), .Q(n2498) );
  OA22X1 U1957 ( .IN1(n3717), .IN2(n3090), .IN3(n3714), .IN4(n3229), .Q(n2499)
         );
  OA221X1 U1958 ( .IN1(n3711), .IN2(n3097), .IN3(n3708), .IN4(n3472), .IN5(
        n2505), .Q(n2497) );
  OA22X1 U1959 ( .IN1(n3705), .IN2(n3089), .IN3(n3702), .IN4(n3228), .Q(n2505)
         );
  OA221X1 U1960 ( .IN1(n3699), .IN2(n3096), .IN3(n3696), .IN4(n3471), .IN5(
        n2507), .Q(n2496) );
  OA22X1 U1961 ( .IN1(n3693), .IN2(n3088), .IN3(n3690), .IN4(n3227), .Q(n2507)
         );
  OA221X1 U1962 ( .IN1(n3687), .IN2(n3095), .IN3(n3684), .IN4(n3470), .IN5(
        n2509), .Q(n2495) );
  OA22X1 U1963 ( .IN1(n3681), .IN2(n3087), .IN3(n3678), .IN4(n3226), .Q(n2509)
         );
  AO22X1 U1964 ( .IN1(n972), .IN2(n3775), .IN3(instr[15]), .IN4(n3765), .Q(
        n932) );
  AO22X1 U1965 ( .IN1(n966), .IN2(n3775), .IN3(instr[14]), .IN4(n3765), .Q(
        n931) );
  AO22X1 U1966 ( .IN1(n973), .IN2(n3775), .IN3(instr[13]), .IN4(n3765), .Q(
        n930) );
  AO22X1 U1967 ( .IN1(n971), .IN2(n3775), .IN3(instr[12]), .IN4(n3765), .Q(
        n929) );
  AO22X1 U1968 ( .IN1(n3814), .IN2(n3775), .IN3(n3767), .IN4(n2511), .Q(n928)
         );
  NAND4X0 U1969 ( .IN1(n2512), .IN2(n2513), .IN3(n2514), .IN4(n2515), .QN(
        n2511) );
  OA221X1 U1970 ( .IN1(n3217), .IN2(n3673), .IN3(n3465), .IN4(n3670), .IN5(
        n2518), .Q(n2515) );
  OA22X1 U1971 ( .IN1(n3086), .IN2(n3667), .IN3(n3345), .IN4(n3664), .Q(n2518)
         );
  OA221X1 U1972 ( .IN1(n3216), .IN2(n3661), .IN3(n3464), .IN4(n3658), .IN5(
        n2523), .Q(n2514) );
  OA22X1 U1973 ( .IN1(n3085), .IN2(n3655), .IN3(n3344), .IN4(n3652), .Q(n2523)
         );
  OA221X1 U1974 ( .IN1(n3215), .IN2(n3649), .IN3(n3463), .IN4(n3646), .IN5(
        n2528), .Q(n2513) );
  OA22X1 U1975 ( .IN1(n3084), .IN2(n3643), .IN3(n3343), .IN4(n3640), .Q(n2528)
         );
  OA221X1 U1976 ( .IN1(n3214), .IN2(n3637), .IN3(n3462), .IN4(n3634), .IN5(
        n2533), .Q(n2512) );
  OA22X1 U1977 ( .IN1(n3083), .IN2(n3631), .IN3(n3342), .IN4(n3628), .Q(n2533)
         );
  AO22X1 U1978 ( .IN1(n3815), .IN2(n3775), .IN3(n3766), .IN4(n2536), .Q(n927)
         );
  NAND4X0 U1979 ( .IN1(n2537), .IN2(n2538), .IN3(n2539), .IN4(n2540), .QN(
        n2536) );
  OA221X1 U1980 ( .IN1(n3213), .IN2(n3673), .IN3(n3461), .IN4(n3670), .IN5(
        n2541), .Q(n2540) );
  OA22X1 U1981 ( .IN1(n3082), .IN2(n3667), .IN3(n3341), .IN4(n3664), .Q(n2541)
         );
  OA221X1 U1982 ( .IN1(n3212), .IN2(n3661), .IN3(n3460), .IN4(n3658), .IN5(
        n2542), .Q(n2539) );
  OA22X1 U1983 ( .IN1(n3081), .IN2(n3655), .IN3(n3340), .IN4(n3652), .Q(n2542)
         );
  OA221X1 U1984 ( .IN1(n3211), .IN2(n3649), .IN3(n3459), .IN4(n3646), .IN5(
        n2543), .Q(n2538) );
  OA22X1 U1985 ( .IN1(n3080), .IN2(n3643), .IN3(n3339), .IN4(n3640), .Q(n2543)
         );
  OA221X1 U1986 ( .IN1(n3210), .IN2(n3637), .IN3(n3458), .IN4(n3634), .IN5(
        n2544), .Q(n2537) );
  OA22X1 U1987 ( .IN1(n3079), .IN2(n3631), .IN3(n3338), .IN4(n3628), .Q(n2544)
         );
  AO22X1 U1988 ( .IN1(n3816), .IN2(n3775), .IN3(n3766), .IN4(n2545), .Q(n926)
         );
  NAND4X0 U1989 ( .IN1(n2546), .IN2(n2547), .IN3(n2548), .IN4(n2549), .QN(
        n2545) );
  OA221X1 U1990 ( .IN1(n3209), .IN2(n3673), .IN3(n3457), .IN4(n3670), .IN5(
        n2550), .Q(n2549) );
  OA22X1 U1991 ( .IN1(n3078), .IN2(n3667), .IN3(n3337), .IN4(n3664), .Q(n2550)
         );
  OA221X1 U1992 ( .IN1(n3208), .IN2(n3661), .IN3(n3456), .IN4(n3658), .IN5(
        n2551), .Q(n2548) );
  OA22X1 U1993 ( .IN1(n3077), .IN2(n3655), .IN3(n3336), .IN4(n3652), .Q(n2551)
         );
  OA221X1 U1994 ( .IN1(n3207), .IN2(n3649), .IN3(n3455), .IN4(n3646), .IN5(
        n2552), .Q(n2547) );
  OA22X1 U1995 ( .IN1(n3076), .IN2(n3643), .IN3(n3335), .IN4(n3640), .Q(n2552)
         );
  OA221X1 U1996 ( .IN1(n3206), .IN2(n3637), .IN3(n3454), .IN4(n3634), .IN5(
        n2553), .Q(n2546) );
  OA22X1 U1997 ( .IN1(n3075), .IN2(n3631), .IN3(n3334), .IN4(n3628), .Q(n2553)
         );
  AO22X1 U1998 ( .IN1(n3817), .IN2(n3775), .IN3(n3766), .IN4(n2554), .Q(n925)
         );
  NAND4X0 U1999 ( .IN1(n2555), .IN2(n2556), .IN3(n2557), .IN4(n2558), .QN(
        n2554) );
  OA221X1 U2000 ( .IN1(n3205), .IN2(n3673), .IN3(n3453), .IN4(n3670), .IN5(
        n2559), .Q(n2558) );
  OA22X1 U2001 ( .IN1(n3074), .IN2(n3667), .IN3(n3333), .IN4(n3664), .Q(n2559)
         );
  OA221X1 U2002 ( .IN1(n3204), .IN2(n3661), .IN3(n3452), .IN4(n3658), .IN5(
        n2560), .Q(n2557) );
  OA22X1 U2003 ( .IN1(n3073), .IN2(n3655), .IN3(n3332), .IN4(n3652), .Q(n2560)
         );
  OA221X1 U2004 ( .IN1(n3203), .IN2(n3649), .IN3(n3451), .IN4(n3646), .IN5(
        n2561), .Q(n2556) );
  OA22X1 U2005 ( .IN1(n3072), .IN2(n3643), .IN3(n3331), .IN4(n3640), .Q(n2561)
         );
  OA221X1 U2006 ( .IN1(n3202), .IN2(n3637), .IN3(n3450), .IN4(n3634), .IN5(
        n2562), .Q(n2555) );
  OA22X1 U2007 ( .IN1(n3071), .IN2(n3631), .IN3(n3330), .IN4(n3628), .Q(n2562)
         );
  AO22X1 U2008 ( .IN1(n3818), .IN2(n3775), .IN3(n3766), .IN4(n2563), .Q(n924)
         );
  NAND4X0 U2009 ( .IN1(n2564), .IN2(n2565), .IN3(n2566), .IN4(n2567), .QN(
        n2563) );
  OA221X1 U2010 ( .IN1(n3201), .IN2(n3673), .IN3(n3449), .IN4(n3670), .IN5(
        n2568), .Q(n2567) );
  OA22X1 U2011 ( .IN1(n3070), .IN2(n3667), .IN3(n3329), .IN4(n3664), .Q(n2568)
         );
  OA221X1 U2012 ( .IN1(n3200), .IN2(n3661), .IN3(n3448), .IN4(n3658), .IN5(
        n2569), .Q(n2566) );
  OA22X1 U2013 ( .IN1(n3069), .IN2(n3655), .IN3(n3328), .IN4(n3652), .Q(n2569)
         );
  OA221X1 U2014 ( .IN1(n3199), .IN2(n3649), .IN3(n3447), .IN4(n3646), .IN5(
        n2570), .Q(n2565) );
  OA22X1 U2015 ( .IN1(n3068), .IN2(n3643), .IN3(n3327), .IN4(n3640), .Q(n2570)
         );
  OA221X1 U2016 ( .IN1(n3198), .IN2(n3637), .IN3(n3446), .IN4(n3634), .IN5(
        n2571), .Q(n2564) );
  OA22X1 U2017 ( .IN1(n3067), .IN2(n3631), .IN3(n3326), .IN4(n3628), .Q(n2571)
         );
  AO22X1 U2018 ( .IN1(n3819), .IN2(n3775), .IN3(n3766), .IN4(n2572), .Q(n923)
         );
  NAND4X0 U2019 ( .IN1(n2573), .IN2(n2574), .IN3(n2575), .IN4(n2576), .QN(
        n2572) );
  OA221X1 U2020 ( .IN1(n3197), .IN2(n3673), .IN3(n3445), .IN4(n3670), .IN5(
        n2577), .Q(n2576) );
  OA22X1 U2021 ( .IN1(n3066), .IN2(n3667), .IN3(n3325), .IN4(n3664), .Q(n2577)
         );
  OA221X1 U2022 ( .IN1(n3196), .IN2(n3661), .IN3(n3444), .IN4(n3658), .IN5(
        n2578), .Q(n2575) );
  OA22X1 U2023 ( .IN1(n3065), .IN2(n3655), .IN3(n3324), .IN4(n3652), .Q(n2578)
         );
  OA221X1 U2024 ( .IN1(n3195), .IN2(n3649), .IN3(n3443), .IN4(n3646), .IN5(
        n2579), .Q(n2574) );
  OA22X1 U2025 ( .IN1(n3064), .IN2(n3643), .IN3(n3323), .IN4(n3640), .Q(n2579)
         );
  OA221X1 U2026 ( .IN1(n3194), .IN2(n3637), .IN3(n3442), .IN4(n3634), .IN5(
        n2580), .Q(n2573) );
  OA22X1 U2027 ( .IN1(n3063), .IN2(n3631), .IN3(n3322), .IN4(n3628), .Q(n2580)
         );
  AO22X1 U2028 ( .IN1(n3820), .IN2(n3775), .IN3(n3766), .IN4(n2581), .Q(n922)
         );
  NAND4X0 U2029 ( .IN1(n2582), .IN2(n2583), .IN3(n2584), .IN4(n2585), .QN(
        n2581) );
  OA221X1 U2030 ( .IN1(n3193), .IN2(n3673), .IN3(n3441), .IN4(n3670), .IN5(
        n2586), .Q(n2585) );
  OA22X1 U2031 ( .IN1(n3062), .IN2(n3667), .IN3(n3321), .IN4(n3664), .Q(n2586)
         );
  OA221X1 U2032 ( .IN1(n3192), .IN2(n3661), .IN3(n3440), .IN4(n3658), .IN5(
        n2587), .Q(n2584) );
  OA22X1 U2033 ( .IN1(n3061), .IN2(n3655), .IN3(n3320), .IN4(n3652), .Q(n2587)
         );
  OA221X1 U2034 ( .IN1(n3191), .IN2(n3649), .IN3(n3439), .IN4(n3646), .IN5(
        n2588), .Q(n2583) );
  OA22X1 U2035 ( .IN1(n3060), .IN2(n3643), .IN3(n3319), .IN4(n3640), .Q(n2588)
         );
  OA221X1 U2036 ( .IN1(n3190), .IN2(n3637), .IN3(n3438), .IN4(n3634), .IN5(
        n2589), .Q(n2582) );
  OA22X1 U2037 ( .IN1(n3059), .IN2(n3631), .IN3(n3318), .IN4(n3628), .Q(n2589)
         );
  AO22X1 U2038 ( .IN1(n3821), .IN2(n3775), .IN3(n3766), .IN4(n2590), .Q(n921)
         );
  NAND4X0 U2039 ( .IN1(n2591), .IN2(n2592), .IN3(n2593), .IN4(n2594), .QN(
        n2590) );
  OA221X1 U2040 ( .IN1(n3189), .IN2(n3673), .IN3(n3437), .IN4(n3670), .IN5(
        n2595), .Q(n2594) );
  OA22X1 U2041 ( .IN1(n3058), .IN2(n3667), .IN3(n3317), .IN4(n3664), .Q(n2595)
         );
  OA221X1 U2042 ( .IN1(n3188), .IN2(n3661), .IN3(n3436), .IN4(n3658), .IN5(
        n2596), .Q(n2593) );
  OA22X1 U2043 ( .IN1(n3057), .IN2(n3655), .IN3(n3316), .IN4(n3652), .Q(n2596)
         );
  OA221X1 U2044 ( .IN1(n3187), .IN2(n3649), .IN3(n3435), .IN4(n3646), .IN5(
        n2597), .Q(n2592) );
  OA22X1 U2045 ( .IN1(n3056), .IN2(n3643), .IN3(n3315), .IN4(n3640), .Q(n2597)
         );
  OA221X1 U2046 ( .IN1(n3186), .IN2(n3637), .IN3(n3434), .IN4(n3634), .IN5(
        n2598), .Q(n2591) );
  OA22X1 U2047 ( .IN1(n3055), .IN2(n3631), .IN3(n3314), .IN4(n3628), .Q(n2598)
         );
  AO22X1 U2048 ( .IN1(n3822), .IN2(n3775), .IN3(n3766), .IN4(n2599), .Q(n920)
         );
  NAND4X0 U2049 ( .IN1(n2600), .IN2(n2601), .IN3(n2602), .IN4(n2603), .QN(
        n2599) );
  OA221X1 U2050 ( .IN1(n3185), .IN2(n3673), .IN3(n3433), .IN4(n3670), .IN5(
        n2604), .Q(n2603) );
  OA22X1 U2051 ( .IN1(n3054), .IN2(n3667), .IN3(n3313), .IN4(n3664), .Q(n2604)
         );
  OA221X1 U2052 ( .IN1(n3184), .IN2(n3661), .IN3(n3432), .IN4(n3658), .IN5(
        n2605), .Q(n2602) );
  OA22X1 U2053 ( .IN1(n3053), .IN2(n3655), .IN3(n3312), .IN4(n3652), .Q(n2605)
         );
  OA221X1 U2054 ( .IN1(n3183), .IN2(n3649), .IN3(n3431), .IN4(n3646), .IN5(
        n2606), .Q(n2601) );
  OA22X1 U2055 ( .IN1(n3052), .IN2(n3643), .IN3(n3311), .IN4(n3640), .Q(n2606)
         );
  OA221X1 U2056 ( .IN1(n3182), .IN2(n3637), .IN3(n3430), .IN4(n3634), .IN5(
        n2607), .Q(n2600) );
  OA22X1 U2057 ( .IN1(n3051), .IN2(n3631), .IN3(n3310), .IN4(n3628), .Q(n2607)
         );
  AO22X1 U2058 ( .IN1(n3823), .IN2(n3775), .IN3(n3766), .IN4(n2608), .Q(n919)
         );
  NAND4X0 U2059 ( .IN1(n2609), .IN2(n2610), .IN3(n2611), .IN4(n2612), .QN(
        n2608) );
  OA221X1 U2060 ( .IN1(n3181), .IN2(n3673), .IN3(n3429), .IN4(n3670), .IN5(
        n2613), .Q(n2612) );
  OA22X1 U2061 ( .IN1(n3050), .IN2(n3667), .IN3(n3309), .IN4(n3664), .Q(n2613)
         );
  OA221X1 U2062 ( .IN1(n3180), .IN2(n3661), .IN3(n3428), .IN4(n3658), .IN5(
        n2614), .Q(n2611) );
  OA22X1 U2063 ( .IN1(n3049), .IN2(n3655), .IN3(n3308), .IN4(n3652), .Q(n2614)
         );
  OA221X1 U2064 ( .IN1(n3179), .IN2(n3649), .IN3(n3427), .IN4(n3646), .IN5(
        n2615), .Q(n2610) );
  OA22X1 U2065 ( .IN1(n3048), .IN2(n3643), .IN3(n3307), .IN4(n3640), .Q(n2615)
         );
  OA221X1 U2066 ( .IN1(n3178), .IN2(n3637), .IN3(n3426), .IN4(n3634), .IN5(
        n2616), .Q(n2609) );
  OA22X1 U2067 ( .IN1(n3047), .IN2(n3631), .IN3(n3306), .IN4(n3628), .Q(n2616)
         );
  AO22X1 U2068 ( .IN1(n3824), .IN2(n3776), .IN3(n3766), .IN4(n2617), .Q(n918)
         );
  NAND4X0 U2069 ( .IN1(n2618), .IN2(n2619), .IN3(n2620), .IN4(n2621), .QN(
        n2617) );
  OA221X1 U2070 ( .IN1(n3177), .IN2(n3673), .IN3(n3425), .IN4(n3670), .IN5(
        n2622), .Q(n2621) );
  OA22X1 U2071 ( .IN1(n3046), .IN2(n3667), .IN3(n3305), .IN4(n3664), .Q(n2622)
         );
  OA221X1 U2072 ( .IN1(n3176), .IN2(n3661), .IN3(n3424), .IN4(n3658), .IN5(
        n2623), .Q(n2620) );
  OA22X1 U2073 ( .IN1(n3045), .IN2(n3655), .IN3(n3304), .IN4(n3652), .Q(n2623)
         );
  OA221X1 U2074 ( .IN1(n3175), .IN2(n3649), .IN3(n3423), .IN4(n3646), .IN5(
        n2624), .Q(n2619) );
  OA22X1 U2075 ( .IN1(n3044), .IN2(n3643), .IN3(n3303), .IN4(n3640), .Q(n2624)
         );
  OA221X1 U2076 ( .IN1(n3174), .IN2(n3637), .IN3(n3422), .IN4(n3634), .IN5(
        n2625), .Q(n2618) );
  OA22X1 U2077 ( .IN1(n3043), .IN2(n3631), .IN3(n3302), .IN4(n3628), .Q(n2625)
         );
  AO22X1 U2078 ( .IN1(n3825), .IN2(n3776), .IN3(n3766), .IN4(n2626), .Q(n917)
         );
  NAND4X0 U2079 ( .IN1(n2627), .IN2(n2628), .IN3(n2629), .IN4(n2630), .QN(
        n2626) );
  OA221X1 U2080 ( .IN1(n3173), .IN2(n3673), .IN3(n3421), .IN4(n3670), .IN5(
        n2631), .Q(n2630) );
  OA22X1 U2081 ( .IN1(n3042), .IN2(n3667), .IN3(n3301), .IN4(n3664), .Q(n2631)
         );
  OA221X1 U2082 ( .IN1(n3172), .IN2(n3661), .IN3(n3420), .IN4(n3658), .IN5(
        n2632), .Q(n2629) );
  OA22X1 U2083 ( .IN1(n3041), .IN2(n3655), .IN3(n3300), .IN4(n3652), .Q(n2632)
         );
  OA221X1 U2084 ( .IN1(n3171), .IN2(n3649), .IN3(n3419), .IN4(n3646), .IN5(
        n2633), .Q(n2628) );
  OA22X1 U2085 ( .IN1(n3040), .IN2(n3643), .IN3(n3299), .IN4(n3640), .Q(n2633)
         );
  OA221X1 U2086 ( .IN1(n3170), .IN2(n3637), .IN3(n3418), .IN4(n3634), .IN5(
        n2634), .Q(n2627) );
  OA22X1 U2087 ( .IN1(n3039), .IN2(n3631), .IN3(n3298), .IN4(n3628), .Q(n2634)
         );
  AO22X1 U2088 ( .IN1(n3826), .IN2(n3776), .IN3(n3766), .IN4(n2635), .Q(n916)
         );
  NAND4X0 U2089 ( .IN1(n2636), .IN2(n2637), .IN3(n2638), .IN4(n2639), .QN(
        n2635) );
  OA221X1 U2090 ( .IN1(n3169), .IN2(n3674), .IN3(n3417), .IN4(n3671), .IN5(
        n2640), .Q(n2639) );
  OA22X1 U2091 ( .IN1(n3038), .IN2(n3668), .IN3(n3297), .IN4(n3665), .Q(n2640)
         );
  OA221X1 U2092 ( .IN1(n3168), .IN2(n3662), .IN3(n3416), .IN4(n3659), .IN5(
        n2641), .Q(n2638) );
  OA22X1 U2093 ( .IN1(n3037), .IN2(n3656), .IN3(n3296), .IN4(n3653), .Q(n2641)
         );
  OA221X1 U2094 ( .IN1(n3167), .IN2(n3650), .IN3(n3415), .IN4(n3647), .IN5(
        n2642), .Q(n2637) );
  OA22X1 U2095 ( .IN1(n3036), .IN2(n3644), .IN3(n3295), .IN4(n3641), .Q(n2642)
         );
  OA221X1 U2096 ( .IN1(n3166), .IN2(n3638), .IN3(n3414), .IN4(n3635), .IN5(
        n2643), .Q(n2636) );
  OA22X1 U2097 ( .IN1(n3035), .IN2(n3632), .IN3(n3294), .IN4(n3629), .Q(n2643)
         );
  AO22X1 U2098 ( .IN1(n3827), .IN2(n3776), .IN3(n3766), .IN4(n2644), .Q(n915)
         );
  NAND4X0 U2099 ( .IN1(n2645), .IN2(n2646), .IN3(n2647), .IN4(n2648), .QN(
        n2644) );
  OA221X1 U2100 ( .IN1(n3165), .IN2(n3674), .IN3(n3413), .IN4(n3671), .IN5(
        n2649), .Q(n2648) );
  OA22X1 U2101 ( .IN1(n3034), .IN2(n3668), .IN3(n3293), .IN4(n3665), .Q(n2649)
         );
  OA221X1 U2102 ( .IN1(n3164), .IN2(n3662), .IN3(n3412), .IN4(n3659), .IN5(
        n2650), .Q(n2647) );
  OA22X1 U2103 ( .IN1(n3033), .IN2(n3656), .IN3(n3292), .IN4(n3653), .Q(n2650)
         );
  OA221X1 U2104 ( .IN1(n3163), .IN2(n3650), .IN3(n3411), .IN4(n3647), .IN5(
        n2651), .Q(n2646) );
  OA22X1 U2105 ( .IN1(n3032), .IN2(n3644), .IN3(n3291), .IN4(n3641), .Q(n2651)
         );
  OA221X1 U2106 ( .IN1(n3162), .IN2(n3638), .IN3(n3410), .IN4(n3635), .IN5(
        n2652), .Q(n2645) );
  OA22X1 U2107 ( .IN1(n3031), .IN2(n3632), .IN3(n3290), .IN4(n3629), .Q(n2652)
         );
  AO22X1 U2108 ( .IN1(n3828), .IN2(n3776), .IN3(n3766), .IN4(n2653), .Q(n914)
         );
  NAND4X0 U2109 ( .IN1(n2654), .IN2(n2655), .IN3(n2656), .IN4(n2657), .QN(
        n2653) );
  OA221X1 U2110 ( .IN1(n3161), .IN2(n3674), .IN3(n3409), .IN4(n3671), .IN5(
        n2658), .Q(n2657) );
  OA22X1 U2111 ( .IN1(n3030), .IN2(n3668), .IN3(n3289), .IN4(n3665), .Q(n2658)
         );
  OA221X1 U2112 ( .IN1(n3160), .IN2(n3662), .IN3(n3408), .IN4(n3659), .IN5(
        n2659), .Q(n2656) );
  OA22X1 U2113 ( .IN1(n3029), .IN2(n3656), .IN3(n3288), .IN4(n3653), .Q(n2659)
         );
  OA221X1 U2114 ( .IN1(n3159), .IN2(n3650), .IN3(n3407), .IN4(n3647), .IN5(
        n2660), .Q(n2655) );
  OA22X1 U2115 ( .IN1(n3028), .IN2(n3644), .IN3(n3287), .IN4(n3641), .Q(n2660)
         );
  OA221X1 U2116 ( .IN1(n3158), .IN2(n3638), .IN3(n3406), .IN4(n3635), .IN5(
        n2661), .Q(n2654) );
  OA22X1 U2117 ( .IN1(n3027), .IN2(n3632), .IN3(n3286), .IN4(n3629), .Q(n2661)
         );
  AO22X1 U2118 ( .IN1(n3829), .IN2(n3776), .IN3(n3766), .IN4(n2662), .Q(n913)
         );
  NAND4X0 U2119 ( .IN1(n2663), .IN2(n2664), .IN3(n2665), .IN4(n2666), .QN(
        n2662) );
  OA221X1 U2120 ( .IN1(n3157), .IN2(n3674), .IN3(n3405), .IN4(n3671), .IN5(
        n2667), .Q(n2666) );
  OA22X1 U2121 ( .IN1(n3026), .IN2(n3668), .IN3(n3285), .IN4(n3665), .Q(n2667)
         );
  OA221X1 U2122 ( .IN1(n3156), .IN2(n3662), .IN3(n3404), .IN4(n3659), .IN5(
        n2668), .Q(n2665) );
  OA22X1 U2123 ( .IN1(n3025), .IN2(n3656), .IN3(n3284), .IN4(n3653), .Q(n2668)
         );
  OA221X1 U2124 ( .IN1(n3155), .IN2(n3650), .IN3(n3403), .IN4(n3647), .IN5(
        n2669), .Q(n2664) );
  OA22X1 U2125 ( .IN1(n3024), .IN2(n3644), .IN3(n3283), .IN4(n3641), .Q(n2669)
         );
  OA221X1 U2126 ( .IN1(n3154), .IN2(n3638), .IN3(n3402), .IN4(n3635), .IN5(
        n2670), .Q(n2663) );
  OA22X1 U2127 ( .IN1(n3023), .IN2(n3632), .IN3(n3282), .IN4(n3629), .Q(n2670)
         );
  AO22X1 U2128 ( .IN1(n3830), .IN2(n3776), .IN3(n3766), .IN4(n2671), .Q(n912)
         );
  NAND4X0 U2129 ( .IN1(n2672), .IN2(n2673), .IN3(n2674), .IN4(n2675), .QN(
        n2671) );
  OA221X1 U2130 ( .IN1(n3153), .IN2(n3674), .IN3(n3401), .IN4(n3671), .IN5(
        n2676), .Q(n2675) );
  OA22X1 U2131 ( .IN1(n3022), .IN2(n3668), .IN3(n3281), .IN4(n3665), .Q(n2676)
         );
  OA221X1 U2132 ( .IN1(n3152), .IN2(n3662), .IN3(n3400), .IN4(n3659), .IN5(
        n2677), .Q(n2674) );
  OA22X1 U2133 ( .IN1(n3021), .IN2(n3656), .IN3(n3280), .IN4(n3653), .Q(n2677)
         );
  OA221X1 U2134 ( .IN1(n3151), .IN2(n3650), .IN3(n3399), .IN4(n3647), .IN5(
        n2678), .Q(n2673) );
  OA22X1 U2135 ( .IN1(n3020), .IN2(n3644), .IN3(n3279), .IN4(n3641), .Q(n2678)
         );
  OA221X1 U2136 ( .IN1(n3150), .IN2(n3638), .IN3(n3398), .IN4(n3635), .IN5(
        n2679), .Q(n2672) );
  OA22X1 U2137 ( .IN1(n3019), .IN2(n3632), .IN3(n3278), .IN4(n3629), .Q(n2679)
         );
  AO22X1 U2138 ( .IN1(n3831), .IN2(n3776), .IN3(n3766), .IN4(n2680), .Q(n911)
         );
  NAND4X0 U2139 ( .IN1(n2681), .IN2(n2682), .IN3(n2683), .IN4(n2684), .QN(
        n2680) );
  OA221X1 U2140 ( .IN1(n3149), .IN2(n3674), .IN3(n3397), .IN4(n3671), .IN5(
        n2685), .Q(n2684) );
  OA22X1 U2141 ( .IN1(n3018), .IN2(n3668), .IN3(n3277), .IN4(n3665), .Q(n2685)
         );
  OA221X1 U2142 ( .IN1(n3148), .IN2(n3662), .IN3(n3396), .IN4(n3659), .IN5(
        n2686), .Q(n2683) );
  OA22X1 U2143 ( .IN1(n3017), .IN2(n3656), .IN3(n3276), .IN4(n3653), .Q(n2686)
         );
  OA221X1 U2144 ( .IN1(n3147), .IN2(n3650), .IN3(n3395), .IN4(n3647), .IN5(
        n2687), .Q(n2682) );
  OA22X1 U2145 ( .IN1(n3016), .IN2(n3644), .IN3(n3275), .IN4(n3641), .Q(n2687)
         );
  OA221X1 U2146 ( .IN1(n3146), .IN2(n3638), .IN3(n3394), .IN4(n3635), .IN5(
        n2688), .Q(n2681) );
  OA22X1 U2147 ( .IN1(n3015), .IN2(n3632), .IN3(n3274), .IN4(n3629), .Q(n2688)
         );
  AO22X1 U2148 ( .IN1(n3832), .IN2(n3776), .IN3(n3766), .IN4(n2689), .Q(n910)
         );
  NAND4X0 U2149 ( .IN1(n2690), .IN2(n2691), .IN3(n2692), .IN4(n2693), .QN(
        n2689) );
  OA221X1 U2150 ( .IN1(n3145), .IN2(n3674), .IN3(n3393), .IN4(n3671), .IN5(
        n2694), .Q(n2693) );
  OA22X1 U2151 ( .IN1(n3014), .IN2(n3668), .IN3(n3273), .IN4(n3665), .Q(n2694)
         );
  OA221X1 U2152 ( .IN1(n3144), .IN2(n3662), .IN3(n3392), .IN4(n3659), .IN5(
        n2695), .Q(n2692) );
  OA22X1 U2153 ( .IN1(n3013), .IN2(n3656), .IN3(n3272), .IN4(n3653), .Q(n2695)
         );
  OA221X1 U2154 ( .IN1(n3143), .IN2(n3650), .IN3(n3391), .IN4(n3647), .IN5(
        n2696), .Q(n2691) );
  OA22X1 U2155 ( .IN1(n3012), .IN2(n3644), .IN3(n3271), .IN4(n3641), .Q(n2696)
         );
  OA221X1 U2156 ( .IN1(n3142), .IN2(n3638), .IN3(n3390), .IN4(n3635), .IN5(
        n2697), .Q(n2690) );
  OA22X1 U2157 ( .IN1(n3011), .IN2(n3632), .IN3(n3270), .IN4(n3629), .Q(n2697)
         );
  AO22X1 U2158 ( .IN1(n3833), .IN2(n3776), .IN3(n3766), .IN4(n2698), .Q(n909)
         );
  NAND4X0 U2159 ( .IN1(n2699), .IN2(n2700), .IN3(n2701), .IN4(n2702), .QN(
        n2698) );
  OA221X1 U2160 ( .IN1(n3141), .IN2(n3674), .IN3(n3389), .IN4(n3671), .IN5(
        n2703), .Q(n2702) );
  OA22X1 U2161 ( .IN1(n3010), .IN2(n3668), .IN3(n3269), .IN4(n3665), .Q(n2703)
         );
  OA221X1 U2162 ( .IN1(n3140), .IN2(n3662), .IN3(n3388), .IN4(n3659), .IN5(
        n2704), .Q(n2701) );
  OA22X1 U2163 ( .IN1(n3009), .IN2(n3656), .IN3(n3268), .IN4(n3653), .Q(n2704)
         );
  OA221X1 U2164 ( .IN1(n3139), .IN2(n3650), .IN3(n3387), .IN4(n3647), .IN5(
        n2705), .Q(n2700) );
  OA22X1 U2165 ( .IN1(n3008), .IN2(n3644), .IN3(n3267), .IN4(n3641), .Q(n2705)
         );
  OA221X1 U2166 ( .IN1(n3138), .IN2(n3638), .IN3(n3386), .IN4(n3635), .IN5(
        n2706), .Q(n2699) );
  OA22X1 U2167 ( .IN1(n3007), .IN2(n3632), .IN3(n3266), .IN4(n3629), .Q(n2706)
         );
  AO22X1 U2168 ( .IN1(n3834), .IN2(n3776), .IN3(n3766), .IN4(n2707), .Q(n908)
         );
  NAND4X0 U2169 ( .IN1(n2708), .IN2(n2709), .IN3(n2710), .IN4(n2711), .QN(
        n2707) );
  OA221X1 U2170 ( .IN1(n3137), .IN2(n3674), .IN3(n3385), .IN4(n3671), .IN5(
        n2712), .Q(n2711) );
  OA22X1 U2171 ( .IN1(n3006), .IN2(n3668), .IN3(n3265), .IN4(n3665), .Q(n2712)
         );
  OA221X1 U2172 ( .IN1(n3136), .IN2(n3662), .IN3(n3384), .IN4(n3659), .IN5(
        n2713), .Q(n2710) );
  OA22X1 U2173 ( .IN1(n3005), .IN2(n3656), .IN3(n3264), .IN4(n3653), .Q(n2713)
         );
  OA221X1 U2174 ( .IN1(n3135), .IN2(n3650), .IN3(n3383), .IN4(n3647), .IN5(
        n2714), .Q(n2709) );
  OA22X1 U2175 ( .IN1(n3004), .IN2(n3644), .IN3(n3263), .IN4(n3641), .Q(n2714)
         );
  OA221X1 U2176 ( .IN1(n3134), .IN2(n3638), .IN3(n3382), .IN4(n3635), .IN5(
        n2715), .Q(n2708) );
  OA22X1 U2177 ( .IN1(n3003), .IN2(n3632), .IN3(n3262), .IN4(n3629), .Q(n2715)
         );
  AO22X1 U2178 ( .IN1(n3835), .IN2(n3776), .IN3(n3766), .IN4(n2716), .Q(n907)
         );
  NAND4X0 U2179 ( .IN1(n2717), .IN2(n2718), .IN3(n2719), .IN4(n2720), .QN(
        n2716) );
  OA221X1 U2180 ( .IN1(n3133), .IN2(n3674), .IN3(n3381), .IN4(n3671), .IN5(
        n2721), .Q(n2720) );
  OA22X1 U2181 ( .IN1(n3002), .IN2(n3668), .IN3(n3261), .IN4(n3665), .Q(n2721)
         );
  OA221X1 U2182 ( .IN1(n3132), .IN2(n3662), .IN3(n3380), .IN4(n3659), .IN5(
        n2722), .Q(n2719) );
  OA22X1 U2183 ( .IN1(n3001), .IN2(n3656), .IN3(n3260), .IN4(n3653), .Q(n2722)
         );
  OA221X1 U2184 ( .IN1(n3131), .IN2(n3650), .IN3(n3379), .IN4(n3647), .IN5(
        n2723), .Q(n2718) );
  OA22X1 U2185 ( .IN1(n3000), .IN2(n3644), .IN3(n3259), .IN4(n3641), .Q(n2723)
         );
  OA221X1 U2186 ( .IN1(n3130), .IN2(n3638), .IN3(n3378), .IN4(n3635), .IN5(
        n2724), .Q(n2717) );
  OA22X1 U2187 ( .IN1(n2999), .IN2(n3632), .IN3(n3258), .IN4(n3629), .Q(n2724)
         );
  AO22X1 U2188 ( .IN1(n3836), .IN2(n3776), .IN3(n3766), .IN4(n2725), .Q(n906)
         );
  NAND4X0 U2189 ( .IN1(n2726), .IN2(n2727), .IN3(n2728), .IN4(n2729), .QN(
        n2725) );
  OA221X1 U2190 ( .IN1(n3129), .IN2(n3674), .IN3(n3377), .IN4(n3671), .IN5(
        n2730), .Q(n2729) );
  OA22X1 U2191 ( .IN1(n2998), .IN2(n3668), .IN3(n3257), .IN4(n3665), .Q(n2730)
         );
  OA221X1 U2192 ( .IN1(n3128), .IN2(n3662), .IN3(n3376), .IN4(n3659), .IN5(
        n2731), .Q(n2728) );
  OA22X1 U2193 ( .IN1(n2997), .IN2(n3656), .IN3(n3256), .IN4(n3653), .Q(n2731)
         );
  OA221X1 U2194 ( .IN1(n3127), .IN2(n3650), .IN3(n3375), .IN4(n3647), .IN5(
        n2732), .Q(n2727) );
  OA22X1 U2195 ( .IN1(n2996), .IN2(n3644), .IN3(n3255), .IN4(n3641), .Q(n2732)
         );
  OA221X1 U2196 ( .IN1(n3126), .IN2(n3638), .IN3(n3374), .IN4(n3635), .IN5(
        n2733), .Q(n2726) );
  OA22X1 U2197 ( .IN1(n2995), .IN2(n3632), .IN3(n3254), .IN4(n3629), .Q(n2733)
         );
  AO22X1 U2198 ( .IN1(n3837), .IN2(n3776), .IN3(n3766), .IN4(n2734), .Q(n905)
         );
  NAND4X0 U2199 ( .IN1(n2735), .IN2(n2736), .IN3(n2737), .IN4(n2738), .QN(
        n2734) );
  OA221X1 U2200 ( .IN1(n3125), .IN2(n3674), .IN3(n3373), .IN4(n3671), .IN5(
        n2739), .Q(n2738) );
  OA22X1 U2201 ( .IN1(n2994), .IN2(n3668), .IN3(n3253), .IN4(n3665), .Q(n2739)
         );
  OA221X1 U2202 ( .IN1(n3124), .IN2(n3662), .IN3(n3372), .IN4(n3659), .IN5(
        n2740), .Q(n2737) );
  OA22X1 U2203 ( .IN1(n2993), .IN2(n3656), .IN3(n3252), .IN4(n3653), .Q(n2740)
         );
  OA221X1 U2204 ( .IN1(n3123), .IN2(n3650), .IN3(n3371), .IN4(n3647), .IN5(
        n2741), .Q(n2736) );
  OA22X1 U2205 ( .IN1(n2992), .IN2(n3644), .IN3(n3251), .IN4(n3641), .Q(n2741)
         );
  OA221X1 U2206 ( .IN1(n3122), .IN2(n3638), .IN3(n3370), .IN4(n3635), .IN5(
        n2742), .Q(n2735) );
  OA22X1 U2207 ( .IN1(n2991), .IN2(n3632), .IN3(n3250), .IN4(n3629), .Q(n2742)
         );
  AO22X1 U2208 ( .IN1(n3838), .IN2(n3777), .IN3(n3766), .IN4(n2743), .Q(n904)
         );
  NAND4X0 U2209 ( .IN1(n2744), .IN2(n2745), .IN3(n2746), .IN4(n2747), .QN(
        n2743) );
  OA221X1 U2210 ( .IN1(n3121), .IN2(n3675), .IN3(n3369), .IN4(n3672), .IN5(
        n2748), .Q(n2747) );
  OA22X1 U2211 ( .IN1(n2990), .IN2(n3669), .IN3(n3249), .IN4(n3666), .Q(n2748)
         );
  OA221X1 U2212 ( .IN1(n3120), .IN2(n3663), .IN3(n3368), .IN4(n3660), .IN5(
        n2749), .Q(n2746) );
  OA22X1 U2213 ( .IN1(n2989), .IN2(n3657), .IN3(n3248), .IN4(n3654), .Q(n2749)
         );
  OA221X1 U2214 ( .IN1(n3119), .IN2(n3651), .IN3(n3367), .IN4(n3648), .IN5(
        n2750), .Q(n2745) );
  OA22X1 U2215 ( .IN1(n2988), .IN2(n3645), .IN3(n3247), .IN4(n3642), .Q(n2750)
         );
  OA221X1 U2216 ( .IN1(n3118), .IN2(n3639), .IN3(n3366), .IN4(n3636), .IN5(
        n2751), .Q(n2744) );
  OA22X1 U2217 ( .IN1(n2987), .IN2(n3633), .IN3(n3246), .IN4(n3630), .Q(n2751)
         );
  AO22X1 U2218 ( .IN1(n3839), .IN2(n3777), .IN3(n3765), .IN4(n2752), .Q(n903)
         );
  NAND4X0 U2219 ( .IN1(n2753), .IN2(n2754), .IN3(n2755), .IN4(n2756), .QN(
        n2752) );
  OA221X1 U2220 ( .IN1(n3117), .IN2(n3675), .IN3(n3365), .IN4(n3672), .IN5(
        n2757), .Q(n2756) );
  OA22X1 U2221 ( .IN1(n2986), .IN2(n3669), .IN3(n3245), .IN4(n3666), .Q(n2757)
         );
  OA221X1 U2222 ( .IN1(n3116), .IN2(n3663), .IN3(n3364), .IN4(n3660), .IN5(
        n2758), .Q(n2755) );
  OA22X1 U2223 ( .IN1(n2985), .IN2(n3657), .IN3(n3244), .IN4(n3654), .Q(n2758)
         );
  OA221X1 U2224 ( .IN1(n3115), .IN2(n3651), .IN3(n3363), .IN4(n3648), .IN5(
        n2759), .Q(n2754) );
  OA22X1 U2225 ( .IN1(n2984), .IN2(n3645), .IN3(n3243), .IN4(n3642), .Q(n2759)
         );
  OA221X1 U2226 ( .IN1(n3114), .IN2(n3639), .IN3(n3362), .IN4(n3636), .IN5(
        n2760), .Q(n2753) );
  OA22X1 U2227 ( .IN1(n2983), .IN2(n3633), .IN3(n3242), .IN4(n3630), .Q(n2760)
         );
  AO22X1 U2228 ( .IN1(n3840), .IN2(n3777), .IN3(n3765), .IN4(n2761), .Q(n902)
         );
  NAND4X0 U2229 ( .IN1(n2762), .IN2(n2763), .IN3(n2764), .IN4(n2765), .QN(
        n2761) );
  OA221X1 U2230 ( .IN1(n3113), .IN2(n3675), .IN3(n3361), .IN4(n3672), .IN5(
        n2766), .Q(n2765) );
  OA22X1 U2231 ( .IN1(n2982), .IN2(n3669), .IN3(n3241), .IN4(n3666), .Q(n2766)
         );
  OA221X1 U2232 ( .IN1(n3112), .IN2(n3663), .IN3(n3360), .IN4(n3660), .IN5(
        n2767), .Q(n2764) );
  OA22X1 U2233 ( .IN1(n2981), .IN2(n3657), .IN3(n3240), .IN4(n3654), .Q(n2767)
         );
  OA221X1 U2234 ( .IN1(n3111), .IN2(n3651), .IN3(n3359), .IN4(n3648), .IN5(
        n2768), .Q(n2763) );
  OA22X1 U2235 ( .IN1(n2980), .IN2(n3645), .IN3(n3239), .IN4(n3642), .Q(n2768)
         );
  OA221X1 U2236 ( .IN1(n3110), .IN2(n3639), .IN3(n3358), .IN4(n3636), .IN5(
        n2769), .Q(n2762) );
  OA22X1 U2237 ( .IN1(n2979), .IN2(n3633), .IN3(n3238), .IN4(n3630), .Q(n2769)
         );
  AO22X1 U2238 ( .IN1(n3841), .IN2(n3777), .IN3(n3765), .IN4(n2770), .Q(n901)
         );
  NAND4X0 U2239 ( .IN1(n2771), .IN2(n2772), .IN3(n2773), .IN4(n2774), .QN(
        n2770) );
  OA221X1 U2240 ( .IN1(n3109), .IN2(n3675), .IN3(n3357), .IN4(n3672), .IN5(
        n2775), .Q(n2774) );
  OA22X1 U2241 ( .IN1(n2978), .IN2(n3669), .IN3(n3237), .IN4(n3666), .Q(n2775)
         );
  OA221X1 U2242 ( .IN1(n3108), .IN2(n3663), .IN3(n3356), .IN4(n3660), .IN5(
        n2776), .Q(n2773) );
  OA22X1 U2243 ( .IN1(n2977), .IN2(n3657), .IN3(n3236), .IN4(n3654), .Q(n2776)
         );
  OA221X1 U2244 ( .IN1(n3107), .IN2(n3651), .IN3(n3355), .IN4(n3648), .IN5(
        n2777), .Q(n2772) );
  OA22X1 U2245 ( .IN1(n2976), .IN2(n3645), .IN3(n3235), .IN4(n3642), .Q(n2777)
         );
  OA221X1 U2246 ( .IN1(n3469), .IN2(n3639), .IN3(n3221), .IN4(n3636), .IN5(
        n2778), .Q(n2771) );
  OA22X1 U2247 ( .IN1(n2975), .IN2(n3633), .IN3(n3234), .IN4(n3630), .Q(n2778)
         );
  AO22X1 U2248 ( .IN1(n3842), .IN2(n3777), .IN3(n3765), .IN4(n2779), .Q(n900)
         );
  NAND4X0 U2249 ( .IN1(n2780), .IN2(n2781), .IN3(n2782), .IN4(n2783), .QN(
        n2779) );
  OA221X1 U2250 ( .IN1(n3106), .IN2(n3675), .IN3(n3354), .IN4(n3672), .IN5(
        n2784), .Q(n2783) );
  OA22X1 U2251 ( .IN1(n2974), .IN2(n3669), .IN3(n3233), .IN4(n3666), .Q(n2784)
         );
  OA221X1 U2252 ( .IN1(n3468), .IN2(n3663), .IN3(n3220), .IN4(n3660), .IN5(
        n2785), .Q(n2782) );
  OA22X1 U2253 ( .IN1(n2973), .IN2(n3657), .IN3(n3232), .IN4(n3654), .Q(n2785)
         );
  OA221X1 U2254 ( .IN1(n3222), .IN2(n3651), .IN3(n3481), .IN4(n3648), .IN5(
        n2786), .Q(n2781) );
  OA22X1 U2255 ( .IN1(n3094), .IN2(n3645), .IN3(n3353), .IN4(n3642), .Q(n2786)
         );
  OA221X1 U2256 ( .IN1(n3105), .IN2(n3639), .IN3(n3480), .IN4(n3636), .IN5(
        n2787), .Q(n2780) );
  OA22X1 U2257 ( .IN1(n3093), .IN2(n3633), .IN3(n3352), .IN4(n3630), .Q(n2787)
         );
  AO22X1 U2258 ( .IN1(n3843), .IN2(n3777), .IN3(n3765), .IN4(n2788), .Q(n899)
         );
  NAND4X0 U2259 ( .IN1(n2789), .IN2(n2790), .IN3(n2791), .IN4(n2792), .QN(
        n2788) );
  OA221X1 U2260 ( .IN1(n3467), .IN2(n3675), .IN3(n3219), .IN4(n3672), .IN5(
        n2793), .Q(n2792) );
  OA22X1 U2261 ( .IN1(n2972), .IN2(n3669), .IN3(n3231), .IN4(n3666), .Q(n2793)
         );
  OA221X1 U2262 ( .IN1(n3104), .IN2(n3663), .IN3(n3479), .IN4(n3660), .IN5(
        n2794), .Q(n2791) );
  OA22X1 U2263 ( .IN1(n3092), .IN2(n3657), .IN3(n3351), .IN4(n3654), .Q(n2794)
         );
  OA221X1 U2264 ( .IN1(n3466), .IN2(n3651), .IN3(n3218), .IN4(n3648), .IN5(
        n2795), .Q(n2790) );
  OA22X1 U2265 ( .IN1(n2971), .IN2(n3645), .IN3(n3230), .IN4(n3642), .Q(n2795)
         );
  OA221X1 U2266 ( .IN1(n3103), .IN2(n3639), .IN3(n3478), .IN4(n3636), .IN5(
        n2796), .Q(n2789) );
  OA22X1 U2267 ( .IN1(n3091), .IN2(n3633), .IN3(n3350), .IN4(n3630), .Q(n2796)
         );
  AO22X1 U2268 ( .IN1(n3844), .IN2(n3777), .IN3(n3767), .IN4(n2797), .Q(n898)
         );
  NAND4X0 U2269 ( .IN1(n2798), .IN2(n2799), .IN3(n2800), .IN4(n2801), .QN(
        n2797) );
  OA221X1 U2270 ( .IN1(n3102), .IN2(n3675), .IN3(n3477), .IN4(n3672), .IN5(
        n2802), .Q(n2801) );
  OA22X1 U2271 ( .IN1(n2970), .IN2(n3669), .IN3(n3349), .IN4(n3666), .Q(n2802)
         );
  OA221X1 U2272 ( .IN1(n3101), .IN2(n3663), .IN3(n3476), .IN4(n3660), .IN5(
        n2803), .Q(n2800) );
  OA22X1 U2273 ( .IN1(n2969), .IN2(n3657), .IN3(n3348), .IN4(n3654), .Q(n2803)
         );
  OA221X1 U2274 ( .IN1(n3100), .IN2(n3651), .IN3(n3475), .IN4(n3648), .IN5(
        n2804), .Q(n2799) );
  OA22X1 U2275 ( .IN1(n2968), .IN2(n3645), .IN3(n3347), .IN4(n3642), .Q(n2804)
         );
  OA221X1 U2276 ( .IN1(n3099), .IN2(n3639), .IN3(n3474), .IN4(n3636), .IN5(
        n2805), .Q(n2798) );
  OA22X1 U2277 ( .IN1(n2967), .IN2(n3633), .IN3(n3346), .IN4(n3630), .Q(n2805)
         );
  AO22X1 U2278 ( .IN1(n3845), .IN2(n3777), .IN3(n3767), .IN4(n2806), .Q(n897)
         );
  NAND4X0 U2279 ( .IN1(n2807), .IN2(n2808), .IN3(n2809), .IN4(n2810), .QN(
        n2806) );
  OA221X1 U2280 ( .IN1(n3098), .IN2(n3675), .IN3(n3473), .IN4(n3672), .IN5(
        n2811), .Q(n2810) );
  OA22X1 U2281 ( .IN1(n3090), .IN2(n3669), .IN3(n3229), .IN4(n3666), .Q(n2811)
         );
  OA221X1 U2282 ( .IN1(n3097), .IN2(n3663), .IN3(n3472), .IN4(n3660), .IN5(
        n2817), .Q(n2809) );
  OA22X1 U2283 ( .IN1(n3089), .IN2(n3657), .IN3(n3228), .IN4(n3654), .Q(n2817)
         );
  OA221X1 U2284 ( .IN1(n3096), .IN2(n3651), .IN3(n3471), .IN4(n3648), .IN5(
        n2819), .Q(n2808) );
  OA22X1 U2285 ( .IN1(n3088), .IN2(n3645), .IN3(n3227), .IN4(n3642), .Q(n2819)
         );
  OA221X1 U2286 ( .IN1(n3095), .IN2(n3639), .IN3(n3470), .IN4(n3636), .IN5(
        n2821), .Q(n2807) );
  OA22X1 U2287 ( .IN1(n3087), .IN2(n3633), .IN3(n3226), .IN4(n3630), .Q(n2821)
         );
  AO22X1 U2288 ( .IN1(IFID_dest[3]), .IN2(n3777), .IN3(instr[3]), .IN4(n3765), 
        .Q(n896) );
  AO22X1 U2289 ( .IN1(IFID_dest[2]), .IN2(n3777), .IN3(instr[2]), .IN4(n3765), 
        .Q(n895) );
  AO22X1 U2290 ( .IN1(IFID_dest[1]), .IN2(n3777), .IN3(instr[1]), .IN4(n3765), 
        .Q(n894) );
  AO22X1 U2291 ( .IN1(IFID_dest[0]), .IN2(n3777), .IN3(instr[0]), .IN4(n3765), 
        .Q(n893) );
  AO22X1 U2292 ( .IN1(\regfile[0][31] ), .IN2(n3624), .IN3(n3625), .IN4(n3778), 
        .Q(n892) );
  AO22X1 U2293 ( .IN1(\regfile[1][31] ), .IN2(n3616), .IN3(n3617), .IN4(n3778), 
        .Q(n891) );
  AO22X1 U2294 ( .IN1(\regfile[2][31] ), .IN2(n3608), .IN3(n3609), .IN4(n3778), 
        .Q(n890) );
  AO22X1 U2295 ( .IN1(\regfile[3][31] ), .IN2(n3600), .IN3(n3601), .IN4(n3778), 
        .Q(n889) );
  AO22X1 U2296 ( .IN1(\regfile[4][31] ), .IN2(n3592), .IN3(n3593), .IN4(n3778), 
        .Q(n888) );
  AO22X1 U2297 ( .IN1(\regfile[5][31] ), .IN2(n3584), .IN3(n3585), .IN4(n3778), 
        .Q(n887) );
  AO22X1 U2298 ( .IN1(\regfile[6][31] ), .IN2(n3576), .IN3(n3577), .IN4(n3778), 
        .Q(n886) );
  AO22X1 U2299 ( .IN1(\regfile[7][31] ), .IN2(n3568), .IN3(n3569), .IN4(n3778), 
        .Q(n885) );
  AO22X1 U2300 ( .IN1(\regfile[8][31] ), .IN2(n3560), .IN3(n3561), .IN4(n3778), 
        .Q(n884) );
  AO22X1 U2301 ( .IN1(\regfile[9][31] ), .IN2(n3552), .IN3(n3553), .IN4(n3778), 
        .Q(n883) );
  AO22X1 U2302 ( .IN1(\regfile[10][31] ), .IN2(n3544), .IN3(n3545), .IN4(n3778), .Q(n882) );
  AO22X1 U2303 ( .IN1(\regfile[11][31] ), .IN2(n3536), .IN3(n3537), .IN4(n3778), .Q(n881) );
  AO22X1 U2304 ( .IN1(\regfile[12][31] ), .IN2(n3528), .IN3(n3529), .IN4(n3778), .Q(n880) );
  AO22X1 U2305 ( .IN1(\regfile[13][31] ), .IN2(n3520), .IN3(n3521), .IN4(n3778), .Q(n879) );
  AO22X1 U2306 ( .IN1(\regfile[14][31] ), .IN2(n3512), .IN3(n3513), .IN4(n3778), .Q(n878) );
  AO22X1 U2307 ( .IN1(\regfile[15][31] ), .IN2(n3504), .IN3(n3505), .IN4(n3778), .Q(n877) );
  AO22X1 U2308 ( .IN1(\regfile[0][30] ), .IN2(n3624), .IN3(n3625), .IN4(n3779), 
        .Q(n876) );
  AO22X1 U2309 ( .IN1(\regfile[1][30] ), .IN2(n3616), .IN3(n3617), .IN4(n3779), 
        .Q(n875) );
  AO22X1 U2310 ( .IN1(\regfile[2][30] ), .IN2(n3608), .IN3(n3609), .IN4(n3779), 
        .Q(n874) );
  AO22X1 U2311 ( .IN1(\regfile[3][30] ), .IN2(n3600), .IN3(n3601), .IN4(n3779), 
        .Q(n873) );
  AO22X1 U2312 ( .IN1(\regfile[4][30] ), .IN2(n3592), .IN3(n3593), .IN4(n3779), 
        .Q(n872) );
  AO22X1 U2313 ( .IN1(\regfile[5][30] ), .IN2(n3584), .IN3(n3585), .IN4(n3779), 
        .Q(n871) );
  AO22X1 U2314 ( .IN1(\regfile[6][30] ), .IN2(n3576), .IN3(n3577), .IN4(n3779), 
        .Q(n870) );
  AO22X1 U2315 ( .IN1(\regfile[7][30] ), .IN2(n3568), .IN3(n3569), .IN4(n3779), 
        .Q(n869) );
  AO22X1 U2316 ( .IN1(\regfile[8][30] ), .IN2(n3560), .IN3(n3561), .IN4(n3779), 
        .Q(n868) );
  AO22X1 U2317 ( .IN1(\regfile[9][30] ), .IN2(n3552), .IN3(n3553), .IN4(n3779), 
        .Q(n867) );
  AO22X1 U2318 ( .IN1(\regfile[10][30] ), .IN2(n3544), .IN3(n3545), .IN4(n3779), .Q(n866) );
  AO22X1 U2319 ( .IN1(\regfile[11][30] ), .IN2(n3536), .IN3(n3537), .IN4(n3779), .Q(n865) );
  AO22X1 U2320 ( .IN1(\regfile[12][30] ), .IN2(n3528), .IN3(n3529), .IN4(n3779), .Q(n864) );
  AO22X1 U2321 ( .IN1(\regfile[13][30] ), .IN2(n3520), .IN3(n3521), .IN4(n3779), .Q(n863) );
  AO22X1 U2322 ( .IN1(\regfile[14][30] ), .IN2(n3512), .IN3(n3513), .IN4(n3779), .Q(n862) );
  AO22X1 U2323 ( .IN1(\regfile[15][30] ), .IN2(n3504), .IN3(n3505), .IN4(n3779), .Q(n861) );
  AO22X1 U2324 ( .IN1(\regfile[0][29] ), .IN2(n3624), .IN3(n3625), .IN4(n3780), 
        .Q(n860) );
  AO22X1 U2325 ( .IN1(\regfile[1][29] ), .IN2(n3616), .IN3(n3617), .IN4(n3780), 
        .Q(n859) );
  AO22X1 U2326 ( .IN1(\regfile[2][29] ), .IN2(n3608), .IN3(n3609), .IN4(n3780), 
        .Q(n858) );
  AO22X1 U2327 ( .IN1(\regfile[3][29] ), .IN2(n3600), .IN3(n3601), .IN4(n3780), 
        .Q(n857) );
  AO22X1 U2328 ( .IN1(\regfile[4][29] ), .IN2(n3592), .IN3(n3593), .IN4(n3780), 
        .Q(n856) );
  AO22X1 U2329 ( .IN1(\regfile[5][29] ), .IN2(n3584), .IN3(n3585), .IN4(n3780), 
        .Q(n855) );
  AO22X1 U2330 ( .IN1(\regfile[6][29] ), .IN2(n3576), .IN3(n3577), .IN4(n3780), 
        .Q(n854) );
  AO22X1 U2331 ( .IN1(\regfile[7][29] ), .IN2(n3568), .IN3(n3569), .IN4(n3780), 
        .Q(n853) );
  AO22X1 U2332 ( .IN1(\regfile[8][29] ), .IN2(n3560), .IN3(n3561), .IN4(n3780), 
        .Q(n852) );
  AO22X1 U2333 ( .IN1(\regfile[9][29] ), .IN2(n3552), .IN3(n3553), .IN4(n3780), 
        .Q(n851) );
  AO22X1 U2334 ( .IN1(\regfile[10][29] ), .IN2(n3544), .IN3(n3545), .IN4(n3780), .Q(n850) );
  AO22X1 U2335 ( .IN1(\regfile[11][29] ), .IN2(n3536), .IN3(n3537), .IN4(n3780), .Q(n849) );
  AO22X1 U2336 ( .IN1(\regfile[12][29] ), .IN2(n3528), .IN3(n3529), .IN4(n3780), .Q(n848) );
  AO22X1 U2337 ( .IN1(\regfile[13][29] ), .IN2(n3520), .IN3(n3521), .IN4(n3780), .Q(n847) );
  AO22X1 U2338 ( .IN1(\regfile[14][29] ), .IN2(n3512), .IN3(n3513), .IN4(n3780), .Q(n846) );
  AO22X1 U2339 ( .IN1(\regfile[15][29] ), .IN2(n3504), .IN3(n3505), .IN4(n3780), .Q(n845) );
  AO22X1 U2340 ( .IN1(\regfile[0][28] ), .IN2(n3624), .IN3(n3625), .IN4(n3781), 
        .Q(n844) );
  AO22X1 U2341 ( .IN1(\regfile[1][28] ), .IN2(n3616), .IN3(n3617), .IN4(n3781), 
        .Q(n843) );
  AO22X1 U2342 ( .IN1(\regfile[2][28] ), .IN2(n3608), .IN3(n3609), .IN4(n3781), 
        .Q(n842) );
  AO22X1 U2343 ( .IN1(\regfile[3][28] ), .IN2(n3600), .IN3(n3601), .IN4(n3781), 
        .Q(n841) );
  AO22X1 U2344 ( .IN1(\regfile[4][28] ), .IN2(n3592), .IN3(n3593), .IN4(n3781), 
        .Q(n840) );
  AO22X1 U2345 ( .IN1(\regfile[5][28] ), .IN2(n3584), .IN3(n3585), .IN4(n3781), 
        .Q(n839) );
  AO22X1 U2346 ( .IN1(\regfile[6][28] ), .IN2(n3576), .IN3(n3577), .IN4(n3781), 
        .Q(n838) );
  AO22X1 U2347 ( .IN1(\regfile[7][28] ), .IN2(n3568), .IN3(n3569), .IN4(n3781), 
        .Q(n837) );
  AO22X1 U2348 ( .IN1(\regfile[8][28] ), .IN2(n3560), .IN3(n3561), .IN4(n3781), 
        .Q(n836) );
  AO22X1 U2349 ( .IN1(\regfile[9][28] ), .IN2(n3552), .IN3(n3553), .IN4(n3781), 
        .Q(n835) );
  AO22X1 U2350 ( .IN1(\regfile[10][28] ), .IN2(n3544), .IN3(n3545), .IN4(n3781), .Q(n834) );
  AO22X1 U2351 ( .IN1(\regfile[11][28] ), .IN2(n3536), .IN3(n3537), .IN4(n3781), .Q(n833) );
  AO22X1 U2352 ( .IN1(\regfile[12][28] ), .IN2(n3528), .IN3(n3529), .IN4(n3781), .Q(n832) );
  AO22X1 U2353 ( .IN1(\regfile[13][28] ), .IN2(n3520), .IN3(n3521), .IN4(n3781), .Q(n831) );
  AO22X1 U2354 ( .IN1(\regfile[14][28] ), .IN2(n3512), .IN3(n3513), .IN4(n3781), .Q(n830) );
  AO22X1 U2355 ( .IN1(\regfile[15][28] ), .IN2(n3504), .IN3(n3505), .IN4(n3781), .Q(n829) );
  AO22X1 U2356 ( .IN1(\regfile[0][27] ), .IN2(n3624), .IN3(n3625), .IN4(n3782), 
        .Q(n828) );
  AO22X1 U2357 ( .IN1(\regfile[1][27] ), .IN2(n3616), .IN3(n3617), .IN4(n3782), 
        .Q(n827) );
  AO22X1 U2358 ( .IN1(\regfile[2][27] ), .IN2(n3608), .IN3(n3609), .IN4(n3782), 
        .Q(n826) );
  AO22X1 U2359 ( .IN1(\regfile[3][27] ), .IN2(n3600), .IN3(n3601), .IN4(n3782), 
        .Q(n825) );
  AO22X1 U2360 ( .IN1(\regfile[4][27] ), .IN2(n3592), .IN3(n3593), .IN4(n3782), 
        .Q(n824) );
  AO22X1 U2361 ( .IN1(\regfile[5][27] ), .IN2(n3584), .IN3(n3585), .IN4(n3782), 
        .Q(n823) );
  AO22X1 U2362 ( .IN1(\regfile[6][27] ), .IN2(n3576), .IN3(n3577), .IN4(n3782), 
        .Q(n822) );
  AO22X1 U2363 ( .IN1(\regfile[7][27] ), .IN2(n3568), .IN3(n3569), .IN4(n3782), 
        .Q(n821) );
  AO22X1 U2364 ( .IN1(\regfile[8][27] ), .IN2(n3560), .IN3(n3561), .IN4(n3782), 
        .Q(n820) );
  AO22X1 U2365 ( .IN1(\regfile[9][27] ), .IN2(n3552), .IN3(n3553), .IN4(n3782), 
        .Q(n819) );
  AO22X1 U2366 ( .IN1(\regfile[10][27] ), .IN2(n3544), .IN3(n3545), .IN4(n3782), .Q(n818) );
  AO22X1 U2367 ( .IN1(\regfile[11][27] ), .IN2(n3536), .IN3(n3537), .IN4(n3782), .Q(n817) );
  AO22X1 U2368 ( .IN1(\regfile[12][27] ), .IN2(n3528), .IN3(n3529), .IN4(n3782), .Q(n816) );
  AO22X1 U2369 ( .IN1(\regfile[13][27] ), .IN2(n3520), .IN3(n3521), .IN4(n3782), .Q(n815) );
  AO22X1 U2370 ( .IN1(\regfile[14][27] ), .IN2(n3512), .IN3(n3513), .IN4(n3782), .Q(n814) );
  AO22X1 U2371 ( .IN1(\regfile[15][27] ), .IN2(n3504), .IN3(n3505), .IN4(n3782), .Q(n813) );
  AO22X1 U2372 ( .IN1(\regfile[0][26] ), .IN2(n3624), .IN3(n3625), .IN4(n3783), 
        .Q(n812) );
  AO22X1 U2373 ( .IN1(\regfile[1][26] ), .IN2(n3616), .IN3(n3617), .IN4(n3783), 
        .Q(n811) );
  AO22X1 U2374 ( .IN1(\regfile[2][26] ), .IN2(n3608), .IN3(n3609), .IN4(n3783), 
        .Q(n810) );
  AO22X1 U2375 ( .IN1(\regfile[3][26] ), .IN2(n3600), .IN3(n3601), .IN4(n3783), 
        .Q(n809) );
  AO22X1 U2376 ( .IN1(\regfile[4][26] ), .IN2(n3592), .IN3(n3593), .IN4(n3783), 
        .Q(n808) );
  AO22X1 U2377 ( .IN1(\regfile[5][26] ), .IN2(n3584), .IN3(n3585), .IN4(n3783), 
        .Q(n807) );
  AO22X1 U2378 ( .IN1(\regfile[6][26] ), .IN2(n3576), .IN3(n3577), .IN4(n3783), 
        .Q(n806) );
  AO22X1 U2379 ( .IN1(\regfile[7][26] ), .IN2(n3568), .IN3(n3569), .IN4(n3783), 
        .Q(n805) );
  AO22X1 U2380 ( .IN1(\regfile[8][26] ), .IN2(n3560), .IN3(n3561), .IN4(n3783), 
        .Q(n804) );
  AO22X1 U2381 ( .IN1(\regfile[9][26] ), .IN2(n3552), .IN3(n3553), .IN4(n3783), 
        .Q(n803) );
  AO22X1 U2382 ( .IN1(\regfile[10][26] ), .IN2(n3544), .IN3(n3545), .IN4(n3783), .Q(n802) );
  AO22X1 U2383 ( .IN1(\regfile[11][26] ), .IN2(n3536), .IN3(n3537), .IN4(n3783), .Q(n801) );
  AO22X1 U2384 ( .IN1(\regfile[12][26] ), .IN2(n3528), .IN3(n3529), .IN4(n3783), .Q(n800) );
  AO22X1 U2385 ( .IN1(\regfile[13][26] ), .IN2(n3520), .IN3(n3521), .IN4(n3783), .Q(n799) );
  AO22X1 U2386 ( .IN1(\regfile[14][26] ), .IN2(n3512), .IN3(n3513), .IN4(n3783), .Q(n798) );
  AO22X1 U2387 ( .IN1(\regfile[15][26] ), .IN2(n3504), .IN3(n3505), .IN4(n3783), .Q(n797) );
  AO22X1 U2388 ( .IN1(\regfile[0][25] ), .IN2(n3624), .IN3(n3625), .IN4(n3784), 
        .Q(n796) );
  AO22X1 U2389 ( .IN1(\regfile[1][25] ), .IN2(n3616), .IN3(n3617), .IN4(n3784), 
        .Q(n795) );
  AO22X1 U2390 ( .IN1(\regfile[2][25] ), .IN2(n3608), .IN3(n3609), .IN4(n3784), 
        .Q(n794) );
  AO22X1 U2391 ( .IN1(\regfile[3][25] ), .IN2(n3600), .IN3(n3601), .IN4(n3784), 
        .Q(n793) );
  AO22X1 U2392 ( .IN1(\regfile[4][25] ), .IN2(n3592), .IN3(n3593), .IN4(n3784), 
        .Q(n792) );
  AO22X1 U2393 ( .IN1(\regfile[5][25] ), .IN2(n3584), .IN3(n3585), .IN4(n3784), 
        .Q(n791) );
  AO22X1 U2394 ( .IN1(\regfile[6][25] ), .IN2(n3576), .IN3(n3577), .IN4(n3784), 
        .Q(n790) );
  AO22X1 U2395 ( .IN1(\regfile[7][25] ), .IN2(n3568), .IN3(n3569), .IN4(n3784), 
        .Q(n789) );
  AO22X1 U2396 ( .IN1(\regfile[8][25] ), .IN2(n3560), .IN3(n3561), .IN4(n3784), 
        .Q(n788) );
  AO22X1 U2397 ( .IN1(\regfile[9][25] ), .IN2(n3552), .IN3(n3553), .IN4(n3784), 
        .Q(n787) );
  AO22X1 U2398 ( .IN1(\regfile[10][25] ), .IN2(n3544), .IN3(n3545), .IN4(n3784), .Q(n786) );
  AO22X1 U2399 ( .IN1(\regfile[11][25] ), .IN2(n3536), .IN3(n3537), .IN4(n3784), .Q(n785) );
  AO22X1 U2400 ( .IN1(\regfile[12][25] ), .IN2(n3528), .IN3(n3529), .IN4(n3784), .Q(n784) );
  AO22X1 U2401 ( .IN1(\regfile[13][25] ), .IN2(n3520), .IN3(n3521), .IN4(n3784), .Q(n783) );
  AO22X1 U2402 ( .IN1(\regfile[14][25] ), .IN2(n3512), .IN3(n3513), .IN4(n3784), .Q(n782) );
  AO22X1 U2403 ( .IN1(\regfile[15][25] ), .IN2(n3504), .IN3(n3505), .IN4(n3784), .Q(n781) );
  AO22X1 U2404 ( .IN1(\regfile[0][24] ), .IN2(n3623), .IN3(n3625), .IN4(n3785), 
        .Q(n780) );
  AO22X1 U2405 ( .IN1(\regfile[1][24] ), .IN2(n3615), .IN3(n3617), .IN4(n3785), 
        .Q(n779) );
  AO22X1 U2406 ( .IN1(\regfile[2][24] ), .IN2(n3607), .IN3(n3609), .IN4(n3785), 
        .Q(n778) );
  AO22X1 U2407 ( .IN1(\regfile[3][24] ), .IN2(n3599), .IN3(n3601), .IN4(n3785), 
        .Q(n777) );
  AO22X1 U2408 ( .IN1(\regfile[4][24] ), .IN2(n3591), .IN3(n3593), .IN4(n3785), 
        .Q(n776) );
  AO22X1 U2409 ( .IN1(\regfile[5][24] ), .IN2(n3583), .IN3(n3585), .IN4(n3785), 
        .Q(n775) );
  AO22X1 U2410 ( .IN1(\regfile[6][24] ), .IN2(n3575), .IN3(n3577), .IN4(n3785), 
        .Q(n774) );
  AO22X1 U2411 ( .IN1(\regfile[7][24] ), .IN2(n3567), .IN3(n3569), .IN4(n3785), 
        .Q(n773) );
  AO22X1 U2412 ( .IN1(\regfile[8][24] ), .IN2(n3559), .IN3(n3561), .IN4(n3785), 
        .Q(n772) );
  AO22X1 U2413 ( .IN1(\regfile[9][24] ), .IN2(n3551), .IN3(n3553), .IN4(n3785), 
        .Q(n771) );
  AO22X1 U2414 ( .IN1(\regfile[10][24] ), .IN2(n3543), .IN3(n3545), .IN4(n3785), .Q(n770) );
  AO22X1 U2415 ( .IN1(\regfile[11][24] ), .IN2(n3535), .IN3(n3537), .IN4(n3785), .Q(n769) );
  AO22X1 U2416 ( .IN1(\regfile[12][24] ), .IN2(n3527), .IN3(n3529), .IN4(n3785), .Q(n768) );
  AO22X1 U2417 ( .IN1(\regfile[13][24] ), .IN2(n3519), .IN3(n3521), .IN4(n3785), .Q(n767) );
  AO22X1 U2418 ( .IN1(\regfile[14][24] ), .IN2(n3511), .IN3(n3513), .IN4(n3785), .Q(n766) );
  AO22X1 U2419 ( .IN1(\regfile[15][24] ), .IN2(n3503), .IN3(n3505), .IN4(n3785), .Q(n765) );
  AO22X1 U2420 ( .IN1(\regfile[0][23] ), .IN2(n3623), .IN3(n3625), .IN4(n3786), 
        .Q(n764) );
  AO22X1 U2421 ( .IN1(\regfile[1][23] ), .IN2(n3615), .IN3(n3617), .IN4(n3786), 
        .Q(n763) );
  AO22X1 U2422 ( .IN1(\regfile[2][23] ), .IN2(n3607), .IN3(n3609), .IN4(n3786), 
        .Q(n762) );
  AO22X1 U2423 ( .IN1(\regfile[3][23] ), .IN2(n3599), .IN3(n3601), .IN4(n3786), 
        .Q(n761) );
  AO22X1 U2424 ( .IN1(\regfile[4][23] ), .IN2(n3591), .IN3(n3593), .IN4(n3786), 
        .Q(n760) );
  AO22X1 U2425 ( .IN1(\regfile[5][23] ), .IN2(n3583), .IN3(n3585), .IN4(n3786), 
        .Q(n759) );
  AO22X1 U2426 ( .IN1(\regfile[6][23] ), .IN2(n3575), .IN3(n3577), .IN4(n3786), 
        .Q(n758) );
  AO22X1 U2427 ( .IN1(\regfile[7][23] ), .IN2(n3567), .IN3(n3569), .IN4(n3786), 
        .Q(n757) );
  AO22X1 U2428 ( .IN1(\regfile[8][23] ), .IN2(n3559), .IN3(n3561), .IN4(n3786), 
        .Q(n756) );
  AO22X1 U2429 ( .IN1(\regfile[9][23] ), .IN2(n3551), .IN3(n3553), .IN4(n3786), 
        .Q(n755) );
  AO22X1 U2430 ( .IN1(\regfile[10][23] ), .IN2(n3543), .IN3(n3545), .IN4(n3786), .Q(n754) );
  AO22X1 U2431 ( .IN1(\regfile[11][23] ), .IN2(n3535), .IN3(n3537), .IN4(n3786), .Q(n753) );
  AO22X1 U2432 ( .IN1(\regfile[12][23] ), .IN2(n3527), .IN3(n3529), .IN4(n3786), .Q(n752) );
  AO22X1 U2433 ( .IN1(\regfile[13][23] ), .IN2(n3519), .IN3(n3521), .IN4(n3786), .Q(n751) );
  AO22X1 U2434 ( .IN1(\regfile[14][23] ), .IN2(n3511), .IN3(n3513), .IN4(n3786), .Q(n750) );
  AO22X1 U2435 ( .IN1(\regfile[15][23] ), .IN2(n3503), .IN3(n3505), .IN4(n3786), .Q(n749) );
  AO22X1 U2436 ( .IN1(\regfile[0][22] ), .IN2(n3623), .IN3(n3625), .IN4(n3787), 
        .Q(n748) );
  AO22X1 U2437 ( .IN1(\regfile[1][22] ), .IN2(n3615), .IN3(n3617), .IN4(n3787), 
        .Q(n747) );
  AO22X1 U2438 ( .IN1(\regfile[2][22] ), .IN2(n3607), .IN3(n3609), .IN4(n3787), 
        .Q(n746) );
  AO22X1 U2439 ( .IN1(\regfile[3][22] ), .IN2(n3599), .IN3(n3601), .IN4(n3787), 
        .Q(n745) );
  AO22X1 U2440 ( .IN1(\regfile[4][22] ), .IN2(n3591), .IN3(n3593), .IN4(n3787), 
        .Q(n744) );
  AO22X1 U2441 ( .IN1(\regfile[5][22] ), .IN2(n3583), .IN3(n3585), .IN4(n3787), 
        .Q(n743) );
  AO22X1 U2442 ( .IN1(\regfile[6][22] ), .IN2(n3575), .IN3(n3577), .IN4(n3787), 
        .Q(n742) );
  AO22X1 U2443 ( .IN1(\regfile[7][22] ), .IN2(n3567), .IN3(n3569), .IN4(n3787), 
        .Q(n741) );
  AO22X1 U2444 ( .IN1(\regfile[8][22] ), .IN2(n3559), .IN3(n3561), .IN4(n3787), 
        .Q(n740) );
  AO22X1 U2445 ( .IN1(\regfile[9][22] ), .IN2(n3551), .IN3(n3553), .IN4(n3787), 
        .Q(n739) );
  AO22X1 U2446 ( .IN1(\regfile[10][22] ), .IN2(n3543), .IN3(n3545), .IN4(n3787), .Q(n738) );
  AO22X1 U2447 ( .IN1(\regfile[11][22] ), .IN2(n3535), .IN3(n3537), .IN4(n3787), .Q(n737) );
  AO22X1 U2448 ( .IN1(\regfile[12][22] ), .IN2(n3527), .IN3(n3529), .IN4(n3787), .Q(n736) );
  AO22X1 U2449 ( .IN1(\regfile[13][22] ), .IN2(n3519), .IN3(n3521), .IN4(n3787), .Q(n735) );
  AO22X1 U2450 ( .IN1(\regfile[14][22] ), .IN2(n3511), .IN3(n3513), .IN4(n3787), .Q(n734) );
  AO22X1 U2451 ( .IN1(\regfile[15][22] ), .IN2(n3503), .IN3(n3505), .IN4(n3787), .Q(n733) );
  AO22X1 U2452 ( .IN1(\regfile[0][21] ), .IN2(n3623), .IN3(n3625), .IN4(n3788), 
        .Q(n732) );
  AO22X1 U2453 ( .IN1(\regfile[1][21] ), .IN2(n3615), .IN3(n3617), .IN4(n3788), 
        .Q(n731) );
  AO22X1 U2454 ( .IN1(\regfile[2][21] ), .IN2(n3607), .IN3(n3609), .IN4(n3788), 
        .Q(n730) );
  AO22X1 U2455 ( .IN1(\regfile[3][21] ), .IN2(n3599), .IN3(n3601), .IN4(n3788), 
        .Q(n729) );
  AO22X1 U2456 ( .IN1(\regfile[4][21] ), .IN2(n3591), .IN3(n3593), .IN4(n3788), 
        .Q(n728) );
  AO22X1 U2457 ( .IN1(\regfile[5][21] ), .IN2(n3583), .IN3(n3585), .IN4(n3788), 
        .Q(n727) );
  AO22X1 U2458 ( .IN1(\regfile[6][21] ), .IN2(n3575), .IN3(n3577), .IN4(n3788), 
        .Q(n726) );
  AO22X1 U2459 ( .IN1(\regfile[7][21] ), .IN2(n3567), .IN3(n3569), .IN4(n3788), 
        .Q(n725) );
  AO22X1 U2460 ( .IN1(\regfile[8][21] ), .IN2(n3559), .IN3(n3561), .IN4(n3788), 
        .Q(n724) );
  AO22X1 U2461 ( .IN1(\regfile[9][21] ), .IN2(n3551), .IN3(n3553), .IN4(n3788), 
        .Q(n723) );
  AO22X1 U2462 ( .IN1(\regfile[10][21] ), .IN2(n3543), .IN3(n3545), .IN4(n3788), .Q(n722) );
  AO22X1 U2463 ( .IN1(\regfile[11][21] ), .IN2(n3535), .IN3(n3537), .IN4(n3788), .Q(n721) );
  AO22X1 U2464 ( .IN1(\regfile[12][21] ), .IN2(n3527), .IN3(n3529), .IN4(n3788), .Q(n720) );
  AO22X1 U2465 ( .IN1(\regfile[13][21] ), .IN2(n3519), .IN3(n3521), .IN4(n3788), .Q(n719) );
  AO22X1 U2466 ( .IN1(\regfile[14][21] ), .IN2(n3511), .IN3(n3513), .IN4(n3788), .Q(n718) );
  AO22X1 U2467 ( .IN1(\regfile[15][21] ), .IN2(n3503), .IN3(n3505), .IN4(n3788), .Q(n717) );
  AO22X1 U2468 ( .IN1(\regfile[0][20] ), .IN2(n3623), .IN3(n3625), .IN4(n3789), 
        .Q(n716) );
  AO22X1 U2469 ( .IN1(\regfile[1][20] ), .IN2(n3615), .IN3(n3617), .IN4(n3789), 
        .Q(n715) );
  AO22X1 U2470 ( .IN1(\regfile[2][20] ), .IN2(n3607), .IN3(n3609), .IN4(n3789), 
        .Q(n714) );
  AO22X1 U2471 ( .IN1(\regfile[3][20] ), .IN2(n3599), .IN3(n3601), .IN4(n3789), 
        .Q(n713) );
  AO22X1 U2472 ( .IN1(\regfile[4][20] ), .IN2(n3591), .IN3(n3593), .IN4(n3789), 
        .Q(n712) );
  AO22X1 U2473 ( .IN1(\regfile[5][20] ), .IN2(n3583), .IN3(n3585), .IN4(n3789), 
        .Q(n711) );
  AO22X1 U2474 ( .IN1(\regfile[6][20] ), .IN2(n3575), .IN3(n3577), .IN4(n3789), 
        .Q(n710) );
  AO22X1 U2475 ( .IN1(\regfile[7][20] ), .IN2(n3567), .IN3(n3569), .IN4(n3789), 
        .Q(n709) );
  AO22X1 U2476 ( .IN1(\regfile[8][20] ), .IN2(n3559), .IN3(n3561), .IN4(n3789), 
        .Q(n708) );
  AO22X1 U2477 ( .IN1(\regfile[9][20] ), .IN2(n3551), .IN3(n3553), .IN4(n3789), 
        .Q(n707) );
  AO22X1 U2478 ( .IN1(\regfile[10][20] ), .IN2(n3543), .IN3(n3545), .IN4(n3789), .Q(n706) );
  AO22X1 U2479 ( .IN1(\regfile[11][20] ), .IN2(n3535), .IN3(n3537), .IN4(n3789), .Q(n705) );
  AO22X1 U2480 ( .IN1(\regfile[12][20] ), .IN2(n3527), .IN3(n3529), .IN4(n3789), .Q(n704) );
  AO22X1 U2481 ( .IN1(\regfile[13][20] ), .IN2(n3519), .IN3(n3521), .IN4(n3789), .Q(n703) );
  AO22X1 U2482 ( .IN1(\regfile[14][20] ), .IN2(n3511), .IN3(n3513), .IN4(n3789), .Q(n702) );
  AO22X1 U2483 ( .IN1(\regfile[15][20] ), .IN2(n3503), .IN3(n3505), .IN4(n3789), .Q(n701) );
  AO22X1 U2484 ( .IN1(\regfile[0][19] ), .IN2(n3623), .IN3(n3626), .IN4(n3790), 
        .Q(n700) );
  AO22X1 U2485 ( .IN1(\regfile[1][19] ), .IN2(n3615), .IN3(n3618), .IN4(n3790), 
        .Q(n699) );
  AO22X1 U2486 ( .IN1(\regfile[2][19] ), .IN2(n3607), .IN3(n3610), .IN4(n3790), 
        .Q(n698) );
  AO22X1 U2487 ( .IN1(\regfile[3][19] ), .IN2(n3599), .IN3(n3602), .IN4(n3790), 
        .Q(n697) );
  AO22X1 U2488 ( .IN1(\regfile[4][19] ), .IN2(n3591), .IN3(n3594), .IN4(n3790), 
        .Q(n696) );
  AO22X1 U2489 ( .IN1(\regfile[5][19] ), .IN2(n3583), .IN3(n3586), .IN4(n3790), 
        .Q(n695) );
  AO22X1 U2490 ( .IN1(\regfile[6][19] ), .IN2(n3575), .IN3(n3578), .IN4(n3790), 
        .Q(n694) );
  AO22X1 U2491 ( .IN1(\regfile[7][19] ), .IN2(n3567), .IN3(n3570), .IN4(n3790), 
        .Q(n693) );
  AO22X1 U2492 ( .IN1(\regfile[8][19] ), .IN2(n3559), .IN3(n3562), .IN4(n3790), 
        .Q(n692) );
  AO22X1 U2493 ( .IN1(\regfile[9][19] ), .IN2(n3551), .IN3(n3554), .IN4(n3790), 
        .Q(n691) );
  AO22X1 U2494 ( .IN1(\regfile[10][19] ), .IN2(n3543), .IN3(n3546), .IN4(n3790), .Q(n690) );
  AO22X1 U2495 ( .IN1(\regfile[11][19] ), .IN2(n3535), .IN3(n3538), .IN4(n3790), .Q(n689) );
  AO22X1 U2496 ( .IN1(\regfile[12][19] ), .IN2(n3527), .IN3(n3530), .IN4(n3790), .Q(n688) );
  AO22X1 U2497 ( .IN1(\regfile[13][19] ), .IN2(n3519), .IN3(n3522), .IN4(n3790), .Q(n687) );
  AO22X1 U2498 ( .IN1(\regfile[14][19] ), .IN2(n3511), .IN3(n3514), .IN4(n3790), .Q(n686) );
  AO22X1 U2499 ( .IN1(\regfile[15][19] ), .IN2(n3503), .IN3(n3506), .IN4(n3790), .Q(n685) );
  AO22X1 U2500 ( .IN1(\regfile[0][18] ), .IN2(n3623), .IN3(n3626), .IN4(n3791), 
        .Q(n684) );
  AO22X1 U2501 ( .IN1(\regfile[1][18] ), .IN2(n3615), .IN3(n3618), .IN4(n3791), 
        .Q(n683) );
  AO22X1 U2502 ( .IN1(\regfile[2][18] ), .IN2(n3607), .IN3(n3610), .IN4(n3791), 
        .Q(n682) );
  AO22X1 U2503 ( .IN1(\regfile[3][18] ), .IN2(n3599), .IN3(n3602), .IN4(n3791), 
        .Q(n681) );
  AO22X1 U2504 ( .IN1(\regfile[4][18] ), .IN2(n3591), .IN3(n3594), .IN4(n3791), 
        .Q(n680) );
  AO22X1 U2505 ( .IN1(\regfile[5][18] ), .IN2(n3583), .IN3(n3586), .IN4(n3791), 
        .Q(n679) );
  AO22X1 U2506 ( .IN1(\regfile[6][18] ), .IN2(n3575), .IN3(n3578), .IN4(n3791), 
        .Q(n678) );
  AO22X1 U2507 ( .IN1(\regfile[7][18] ), .IN2(n3567), .IN3(n3570), .IN4(n3791), 
        .Q(n677) );
  AO22X1 U2508 ( .IN1(\regfile[8][18] ), .IN2(n3559), .IN3(n3562), .IN4(n3791), 
        .Q(n676) );
  AO22X1 U2509 ( .IN1(\regfile[9][18] ), .IN2(n3551), .IN3(n3554), .IN4(n3791), 
        .Q(n675) );
  AO22X1 U2510 ( .IN1(\regfile[10][18] ), .IN2(n3543), .IN3(n3546), .IN4(n3791), .Q(n674) );
  AO22X1 U2511 ( .IN1(\regfile[11][18] ), .IN2(n3535), .IN3(n3538), .IN4(n3791), .Q(n673) );
  AO22X1 U2512 ( .IN1(\regfile[12][18] ), .IN2(n3527), .IN3(n3530), .IN4(n3791), .Q(n672) );
  AO22X1 U2513 ( .IN1(\regfile[13][18] ), .IN2(n3519), .IN3(n3522), .IN4(n3791), .Q(n671) );
  AO22X1 U2514 ( .IN1(\regfile[14][18] ), .IN2(n3511), .IN3(n3514), .IN4(n3791), .Q(n670) );
  AO22X1 U2515 ( .IN1(\regfile[15][18] ), .IN2(n3503), .IN3(n3506), .IN4(n3791), .Q(n669) );
  AO22X1 U2516 ( .IN1(\regfile[0][17] ), .IN2(n3622), .IN3(n3626), .IN4(n3792), 
        .Q(n668) );
  AO22X1 U2517 ( .IN1(\regfile[1][17] ), .IN2(n3614), .IN3(n3618), .IN4(n3792), 
        .Q(n667) );
  AO22X1 U2518 ( .IN1(\regfile[2][17] ), .IN2(n3606), .IN3(n3610), .IN4(n3792), 
        .Q(n666) );
  AO22X1 U2519 ( .IN1(\regfile[3][17] ), .IN2(n3598), .IN3(n3602), .IN4(n3792), 
        .Q(n665) );
  AO22X1 U2520 ( .IN1(\regfile[4][17] ), .IN2(n3590), .IN3(n3594), .IN4(n3792), 
        .Q(n664) );
  AO22X1 U2521 ( .IN1(\regfile[5][17] ), .IN2(n3582), .IN3(n3586), .IN4(n3792), 
        .Q(n663) );
  AO22X1 U2522 ( .IN1(\regfile[6][17] ), .IN2(n3574), .IN3(n3578), .IN4(n3792), 
        .Q(n662) );
  AO22X1 U2523 ( .IN1(\regfile[7][17] ), .IN2(n3566), .IN3(n3570), .IN4(n3792), 
        .Q(n661) );
  AO22X1 U2524 ( .IN1(\regfile[8][17] ), .IN2(n3558), .IN3(n3562), .IN4(n3792), 
        .Q(n660) );
  AO22X1 U2525 ( .IN1(\regfile[9][17] ), .IN2(n3550), .IN3(n3554), .IN4(n3792), 
        .Q(n659) );
  AO22X1 U2526 ( .IN1(\regfile[10][17] ), .IN2(n3542), .IN3(n3546), .IN4(n3792), .Q(n658) );
  AO22X1 U2527 ( .IN1(\regfile[11][17] ), .IN2(n3534), .IN3(n3538), .IN4(n3792), .Q(n657) );
  AO22X1 U2528 ( .IN1(\regfile[12][17] ), .IN2(n3526), .IN3(n3530), .IN4(n3792), .Q(n656) );
  AO22X1 U2529 ( .IN1(\regfile[13][17] ), .IN2(n3518), .IN3(n3522), .IN4(n3792), .Q(n655) );
  AO22X1 U2530 ( .IN1(\regfile[14][17] ), .IN2(n3510), .IN3(n3514), .IN4(n3792), .Q(n654) );
  AO22X1 U2531 ( .IN1(\regfile[15][17] ), .IN2(n3502), .IN3(n3506), .IN4(n3792), .Q(n653) );
  AO22X1 U2532 ( .IN1(\regfile[0][16] ), .IN2(n3622), .IN3(n3626), .IN4(n3793), 
        .Q(n652) );
  AO22X1 U2533 ( .IN1(\regfile[1][16] ), .IN2(n3614), .IN3(n3618), .IN4(n3793), 
        .Q(n651) );
  AO22X1 U2534 ( .IN1(\regfile[2][16] ), .IN2(n3606), .IN3(n3610), .IN4(n3793), 
        .Q(n650) );
  AO22X1 U2535 ( .IN1(\regfile[3][16] ), .IN2(n3598), .IN3(n3602), .IN4(n3793), 
        .Q(n649) );
  AO22X1 U2536 ( .IN1(\regfile[4][16] ), .IN2(n3590), .IN3(n3594), .IN4(n3793), 
        .Q(n648) );
  AO22X1 U2537 ( .IN1(\regfile[5][16] ), .IN2(n3582), .IN3(n3586), .IN4(n3793), 
        .Q(n647) );
  AO22X1 U2538 ( .IN1(\regfile[6][16] ), .IN2(n3574), .IN3(n3578), .IN4(n3793), 
        .Q(n646) );
  AO22X1 U2539 ( .IN1(\regfile[7][16] ), .IN2(n3566), .IN3(n3570), .IN4(n3793), 
        .Q(n645) );
  AO22X1 U2540 ( .IN1(\regfile[8][16] ), .IN2(n3558), .IN3(n3562), .IN4(n3793), 
        .Q(n644) );
  AO22X1 U2541 ( .IN1(\regfile[9][16] ), .IN2(n3550), .IN3(n3554), .IN4(n3793), 
        .Q(n643) );
  AO22X1 U2542 ( .IN1(\regfile[10][16] ), .IN2(n3542), .IN3(n3546), .IN4(n3793), .Q(n642) );
  AO22X1 U2543 ( .IN1(\regfile[11][16] ), .IN2(n3534), .IN3(n3538), .IN4(n3793), .Q(n641) );
  AO22X1 U2544 ( .IN1(\regfile[12][16] ), .IN2(n3526), .IN3(n3530), .IN4(n3793), .Q(n640) );
  AO22X1 U2545 ( .IN1(\regfile[13][16] ), .IN2(n3518), .IN3(n3522), .IN4(n3793), .Q(n639) );
  AO22X1 U2546 ( .IN1(\regfile[14][16] ), .IN2(n3510), .IN3(n3514), .IN4(n3793), .Q(n638) );
  AO22X1 U2547 ( .IN1(\regfile[15][16] ), .IN2(n3502), .IN3(n3506), .IN4(n3793), .Q(n637) );
  AO22X1 U2548 ( .IN1(\regfile[0][15] ), .IN2(n3622), .IN3(n3626), .IN4(n3794), 
        .Q(n636) );
  AO22X1 U2549 ( .IN1(\regfile[1][15] ), .IN2(n3614), .IN3(n3618), .IN4(n3794), 
        .Q(n635) );
  AO22X1 U2550 ( .IN1(\regfile[2][15] ), .IN2(n3606), .IN3(n3610), .IN4(n3794), 
        .Q(n634) );
  AO22X1 U2551 ( .IN1(\regfile[3][15] ), .IN2(n3598), .IN3(n3602), .IN4(n3794), 
        .Q(n633) );
  AO22X1 U2552 ( .IN1(\regfile[4][15] ), .IN2(n3590), .IN3(n3594), .IN4(n3794), 
        .Q(n632) );
  AO22X1 U2553 ( .IN1(\regfile[5][15] ), .IN2(n3582), .IN3(n3586), .IN4(n3794), 
        .Q(n631) );
  AO22X1 U2554 ( .IN1(\regfile[6][15] ), .IN2(n3574), .IN3(n3578), .IN4(n3794), 
        .Q(n630) );
  AO22X1 U2555 ( .IN1(\regfile[7][15] ), .IN2(n3566), .IN3(n3570), .IN4(n3794), 
        .Q(n629) );
  AO22X1 U2556 ( .IN1(\regfile[8][15] ), .IN2(n3558), .IN3(n3562), .IN4(n3794), 
        .Q(n628) );
  AO22X1 U2557 ( .IN1(\regfile[9][15] ), .IN2(n3550), .IN3(n3554), .IN4(n3794), 
        .Q(n627) );
  AO22X1 U2558 ( .IN1(\regfile[10][15] ), .IN2(n3542), .IN3(n3546), .IN4(n3794), .Q(n626) );
  AO22X1 U2559 ( .IN1(\regfile[11][15] ), .IN2(n3534), .IN3(n3538), .IN4(n3794), .Q(n625) );
  AO22X1 U2560 ( .IN1(\regfile[12][15] ), .IN2(n3526), .IN3(n3530), .IN4(n3794), .Q(n624) );
  AO22X1 U2561 ( .IN1(\regfile[13][15] ), .IN2(n3518), .IN3(n3522), .IN4(n3794), .Q(n623) );
  AO22X1 U2562 ( .IN1(\regfile[14][15] ), .IN2(n3510), .IN3(n3514), .IN4(n3794), .Q(n622) );
  AO22X1 U2563 ( .IN1(\regfile[15][15] ), .IN2(n3502), .IN3(n3506), .IN4(n3794), .Q(n621) );
  AO22X1 U2564 ( .IN1(\regfile[0][14] ), .IN2(n3622), .IN3(n3626), .IN4(n3795), 
        .Q(n620) );
  AO22X1 U2565 ( .IN1(\regfile[1][14] ), .IN2(n3614), .IN3(n3618), .IN4(n3795), 
        .Q(n619) );
  AO22X1 U2566 ( .IN1(\regfile[2][14] ), .IN2(n3606), .IN3(n3610), .IN4(n3795), 
        .Q(n618) );
  AO22X1 U2567 ( .IN1(\regfile[3][14] ), .IN2(n3598), .IN3(n3602), .IN4(n3795), 
        .Q(n617) );
  AO22X1 U2568 ( .IN1(\regfile[4][14] ), .IN2(n3590), .IN3(n3594), .IN4(n3795), 
        .Q(n616) );
  AO22X1 U2569 ( .IN1(\regfile[5][14] ), .IN2(n3582), .IN3(n3586), .IN4(n3795), 
        .Q(n615) );
  AO22X1 U2570 ( .IN1(\regfile[6][14] ), .IN2(n3574), .IN3(n3578), .IN4(n3795), 
        .Q(n614) );
  AO22X1 U2571 ( .IN1(\regfile[7][14] ), .IN2(n3566), .IN3(n3570), .IN4(n3795), 
        .Q(n613) );
  AO22X1 U2572 ( .IN1(\regfile[8][14] ), .IN2(n3558), .IN3(n3562), .IN4(n3795), 
        .Q(n612) );
  AO22X1 U2573 ( .IN1(\regfile[9][14] ), .IN2(n3550), .IN3(n3554), .IN4(n3795), 
        .Q(n611) );
  AO22X1 U2574 ( .IN1(\regfile[10][14] ), .IN2(n3542), .IN3(n3546), .IN4(n3795), .Q(n610) );
  AO22X1 U2575 ( .IN1(\regfile[11][14] ), .IN2(n3534), .IN3(n3538), .IN4(n3795), .Q(n609) );
  AO22X1 U2576 ( .IN1(\regfile[12][14] ), .IN2(n3526), .IN3(n3530), .IN4(n3795), .Q(n608) );
  AO22X1 U2577 ( .IN1(\regfile[13][14] ), .IN2(n3518), .IN3(n3522), .IN4(n3795), .Q(n607) );
  AO22X1 U2578 ( .IN1(\regfile[14][14] ), .IN2(n3510), .IN3(n3514), .IN4(n3795), .Q(n606) );
  AO22X1 U2579 ( .IN1(\regfile[15][14] ), .IN2(n3502), .IN3(n3506), .IN4(n3795), .Q(n605) );
  AO22X1 U2580 ( .IN1(\regfile[0][13] ), .IN2(n3622), .IN3(n3626), .IN4(n3796), 
        .Q(n604) );
  AO22X1 U2581 ( .IN1(\regfile[1][13] ), .IN2(n3614), .IN3(n3618), .IN4(n3796), 
        .Q(n603) );
  AO22X1 U2582 ( .IN1(\regfile[2][13] ), .IN2(n3606), .IN3(n3610), .IN4(n3796), 
        .Q(n602) );
  AO22X1 U2583 ( .IN1(\regfile[3][13] ), .IN2(n3598), .IN3(n3602), .IN4(n3796), 
        .Q(n601) );
  AO22X1 U2584 ( .IN1(\regfile[4][13] ), .IN2(n3590), .IN3(n3594), .IN4(n3796), 
        .Q(n600) );
  AO22X1 U2585 ( .IN1(\regfile[5][13] ), .IN2(n3582), .IN3(n3586), .IN4(n3796), 
        .Q(n599) );
  AO22X1 U2586 ( .IN1(\regfile[6][13] ), .IN2(n3574), .IN3(n3578), .IN4(n3796), 
        .Q(n598) );
  AO22X1 U2587 ( .IN1(\regfile[7][13] ), .IN2(n3566), .IN3(n3570), .IN4(n3796), 
        .Q(n597) );
  AO22X1 U2588 ( .IN1(\regfile[8][13] ), .IN2(n3558), .IN3(n3562), .IN4(n3796), 
        .Q(n596) );
  AO22X1 U2589 ( .IN1(\regfile[9][13] ), .IN2(n3550), .IN3(n3554), .IN4(n3796), 
        .Q(n595) );
  AO22X1 U2590 ( .IN1(\regfile[10][13] ), .IN2(n3542), .IN3(n3546), .IN4(n3796), .Q(n594) );
  AO22X1 U2591 ( .IN1(\regfile[11][13] ), .IN2(n3534), .IN3(n3538), .IN4(n3796), .Q(n593) );
  AO22X1 U2592 ( .IN1(\regfile[12][13] ), .IN2(n3526), .IN3(n3530), .IN4(n3796), .Q(n592) );
  AO22X1 U2593 ( .IN1(\regfile[13][13] ), .IN2(n3518), .IN3(n3522), .IN4(n3796), .Q(n591) );
  AO22X1 U2594 ( .IN1(\regfile[14][13] ), .IN2(n3510), .IN3(n3514), .IN4(n3796), .Q(n590) );
  AO22X1 U2595 ( .IN1(\regfile[15][13] ), .IN2(n3502), .IN3(n3506), .IN4(n3796), .Q(n589) );
  AO22X1 U2596 ( .IN1(\regfile[0][12] ), .IN2(n3622), .IN3(n3626), .IN4(n3797), 
        .Q(n588) );
  AO22X1 U2597 ( .IN1(\regfile[1][12] ), .IN2(n3614), .IN3(n3618), .IN4(n3797), 
        .Q(n587) );
  AO22X1 U2598 ( .IN1(\regfile[2][12] ), .IN2(n3606), .IN3(n3610), .IN4(n3797), 
        .Q(n586) );
  AO22X1 U2599 ( .IN1(\regfile[3][12] ), .IN2(n3598), .IN3(n3602), .IN4(n3797), 
        .Q(n585) );
  AO22X1 U2600 ( .IN1(\regfile[4][12] ), .IN2(n3590), .IN3(n3594), .IN4(n3797), 
        .Q(n584) );
  AO22X1 U2601 ( .IN1(\regfile[5][12] ), .IN2(n3582), .IN3(n3586), .IN4(n3797), 
        .Q(n583) );
  AO22X1 U2602 ( .IN1(\regfile[6][12] ), .IN2(n3574), .IN3(n3578), .IN4(n3797), 
        .Q(n582) );
  AO22X1 U2603 ( .IN1(\regfile[7][12] ), .IN2(n3566), .IN3(n3570), .IN4(n3797), 
        .Q(n581) );
  AO22X1 U2604 ( .IN1(\regfile[8][12] ), .IN2(n3558), .IN3(n3562), .IN4(n3797), 
        .Q(n580) );
  AO22X1 U2605 ( .IN1(\regfile[9][12] ), .IN2(n3550), .IN3(n3554), .IN4(n3797), 
        .Q(n579) );
  AO22X1 U2606 ( .IN1(\regfile[10][12] ), .IN2(n3542), .IN3(n3546), .IN4(n3797), .Q(n578) );
  AO22X1 U2607 ( .IN1(\regfile[11][12] ), .IN2(n3534), .IN3(n3538), .IN4(n3797), .Q(n577) );
  AO22X1 U2608 ( .IN1(\regfile[12][12] ), .IN2(n3526), .IN3(n3530), .IN4(n3797), .Q(n576) );
  AO22X1 U2609 ( .IN1(\regfile[13][12] ), .IN2(n3518), .IN3(n3522), .IN4(n3797), .Q(n575) );
  AO22X1 U2610 ( .IN1(\regfile[14][12] ), .IN2(n3510), .IN3(n3514), .IN4(n3797), .Q(n574) );
  AO22X1 U2611 ( .IN1(\regfile[15][12] ), .IN2(n3502), .IN3(n3506), .IN4(n3797), .Q(n573) );
  AO22X1 U2612 ( .IN1(\regfile[0][11] ), .IN2(n3622), .IN3(n3626), .IN4(n3798), 
        .Q(n572) );
  AO22X1 U2613 ( .IN1(\regfile[1][11] ), .IN2(n3614), .IN3(n3618), .IN4(n3798), 
        .Q(n571) );
  AO22X1 U2614 ( .IN1(\regfile[2][11] ), .IN2(n3606), .IN3(n3610), .IN4(n3798), 
        .Q(n570) );
  AO22X1 U2615 ( .IN1(\regfile[3][11] ), .IN2(n3598), .IN3(n3602), .IN4(n3798), 
        .Q(n569) );
  AO22X1 U2616 ( .IN1(\regfile[4][11] ), .IN2(n3590), .IN3(n3594), .IN4(n3798), 
        .Q(n568) );
  AO22X1 U2617 ( .IN1(\regfile[5][11] ), .IN2(n3582), .IN3(n3586), .IN4(n3798), 
        .Q(n567) );
  AO22X1 U2618 ( .IN1(\regfile[6][11] ), .IN2(n3574), .IN3(n3578), .IN4(n3798), 
        .Q(n566) );
  AO22X1 U2619 ( .IN1(\regfile[7][11] ), .IN2(n3566), .IN3(n3570), .IN4(n3798), 
        .Q(n565) );
  AO22X1 U2620 ( .IN1(\regfile[8][11] ), .IN2(n3558), .IN3(n3562), .IN4(n3798), 
        .Q(n564) );
  AO22X1 U2621 ( .IN1(\regfile[9][11] ), .IN2(n3550), .IN3(n3554), .IN4(n3798), 
        .Q(n563) );
  AO22X1 U2622 ( .IN1(\regfile[10][11] ), .IN2(n3542), .IN3(n3546), .IN4(n3798), .Q(n562) );
  AO22X1 U2623 ( .IN1(\regfile[11][11] ), .IN2(n3534), .IN3(n3538), .IN4(n3798), .Q(n561) );
  AO22X1 U2624 ( .IN1(\regfile[12][11] ), .IN2(n3526), .IN3(n3530), .IN4(n3798), .Q(n560) );
  AO22X1 U2625 ( .IN1(\regfile[13][11] ), .IN2(n3518), .IN3(n3522), .IN4(n3798), .Q(n559) );
  AO22X1 U2626 ( .IN1(\regfile[14][11] ), .IN2(n3510), .IN3(n3514), .IN4(n3798), .Q(n558) );
  AO22X1 U2627 ( .IN1(\regfile[15][11] ), .IN2(n3502), .IN3(n3506), .IN4(n3798), .Q(n557) );
  AO22X1 U2628 ( .IN1(\regfile[0][10] ), .IN2(n3621), .IN3(n3626), .IN4(n3799), 
        .Q(n556) );
  AO22X1 U2629 ( .IN1(\regfile[1][10] ), .IN2(n3613), .IN3(n3618), .IN4(n3799), 
        .Q(n555) );
  AO22X1 U2630 ( .IN1(\regfile[2][10] ), .IN2(n3605), .IN3(n3610), .IN4(n3799), 
        .Q(n554) );
  AO22X1 U2631 ( .IN1(\regfile[3][10] ), .IN2(n3597), .IN3(n3602), .IN4(n3799), 
        .Q(n553) );
  AO22X1 U2632 ( .IN1(\regfile[4][10] ), .IN2(n3589), .IN3(n3594), .IN4(n3799), 
        .Q(n552) );
  AO22X1 U2633 ( .IN1(\regfile[5][10] ), .IN2(n3581), .IN3(n3586), .IN4(n3799), 
        .Q(n551) );
  AO22X1 U2634 ( .IN1(\regfile[6][10] ), .IN2(n3573), .IN3(n3578), .IN4(n3799), 
        .Q(n550) );
  AO22X1 U2635 ( .IN1(\regfile[7][10] ), .IN2(n3565), .IN3(n3570), .IN4(n3799), 
        .Q(n549) );
  AO22X1 U2636 ( .IN1(\regfile[8][10] ), .IN2(n3557), .IN3(n3562), .IN4(n3799), 
        .Q(n548) );
  AO22X1 U2637 ( .IN1(\regfile[9][10] ), .IN2(n3549), .IN3(n3554), .IN4(n3799), 
        .Q(n547) );
  AO22X1 U2638 ( .IN1(\regfile[10][10] ), .IN2(n3541), .IN3(n3546), .IN4(n3799), .Q(n546) );
  AO22X1 U2639 ( .IN1(\regfile[11][10] ), .IN2(n3533), .IN3(n3538), .IN4(n3799), .Q(n545) );
  AO22X1 U2640 ( .IN1(\regfile[12][10] ), .IN2(n3525), .IN3(n3530), .IN4(n3799), .Q(n544) );
  AO22X1 U2641 ( .IN1(\regfile[13][10] ), .IN2(n3517), .IN3(n3522), .IN4(n3799), .Q(n543) );
  AO22X1 U2642 ( .IN1(\regfile[14][10] ), .IN2(n3509), .IN3(n3514), .IN4(n3799), .Q(n542) );
  AO22X1 U2643 ( .IN1(\regfile[15][10] ), .IN2(n3501), .IN3(n3506), .IN4(n3799), .Q(n541) );
  AO22X1 U2644 ( .IN1(\regfile[0][9] ), .IN2(n3621), .IN3(n3626), .IN4(n3800), 
        .Q(n540) );
  AO22X1 U2645 ( .IN1(\regfile[1][9] ), .IN2(n3613), .IN3(n3618), .IN4(n3800), 
        .Q(n539) );
  AO22X1 U2646 ( .IN1(\regfile[2][9] ), .IN2(n3605), .IN3(n3610), .IN4(n3800), 
        .Q(n538) );
  AO22X1 U2647 ( .IN1(\regfile[3][9] ), .IN2(n3597), .IN3(n3602), .IN4(n3800), 
        .Q(n537) );
  AO22X1 U2648 ( .IN1(\regfile[4][9] ), .IN2(n3589), .IN3(n3594), .IN4(n3800), 
        .Q(n536) );
  AO22X1 U2649 ( .IN1(\regfile[5][9] ), .IN2(n3581), .IN3(n3586), .IN4(n3800), 
        .Q(n535) );
  AO22X1 U2650 ( .IN1(\regfile[6][9] ), .IN2(n3573), .IN3(n3578), .IN4(n3800), 
        .Q(n534) );
  AO22X1 U2651 ( .IN1(\regfile[7][9] ), .IN2(n3565), .IN3(n3570), .IN4(n3800), 
        .Q(n533) );
  AO22X1 U2652 ( .IN1(\regfile[8][9] ), .IN2(n3557), .IN3(n3562), .IN4(n3800), 
        .Q(n532) );
  AO22X1 U2653 ( .IN1(\regfile[9][9] ), .IN2(n3549), .IN3(n3554), .IN4(n3800), 
        .Q(n531) );
  AO22X1 U2654 ( .IN1(\regfile[10][9] ), .IN2(n3541), .IN3(n3546), .IN4(n3800), 
        .Q(n530) );
  AO22X1 U2655 ( .IN1(\regfile[11][9] ), .IN2(n3533), .IN3(n3538), .IN4(n3800), 
        .Q(n529) );
  AO22X1 U2656 ( .IN1(\regfile[12][9] ), .IN2(n3525), .IN3(n3530), .IN4(n3800), 
        .Q(n528) );
  AO22X1 U2657 ( .IN1(\regfile[13][9] ), .IN2(n3517), .IN3(n3522), .IN4(n3800), 
        .Q(n527) );
  AO22X1 U2658 ( .IN1(\regfile[14][9] ), .IN2(n3509), .IN3(n3514), .IN4(n3800), 
        .Q(n526) );
  AO22X1 U2659 ( .IN1(\regfile[15][9] ), .IN2(n3501), .IN3(n3506), .IN4(n3800), 
        .Q(n525) );
  AO22X1 U2660 ( .IN1(\regfile[0][8] ), .IN2(n3621), .IN3(n3626), .IN4(n3801), 
        .Q(n524) );
  AO22X1 U2661 ( .IN1(\regfile[1][8] ), .IN2(n3613), .IN3(n3618), .IN4(n3801), 
        .Q(n523) );
  AO22X1 U2662 ( .IN1(\regfile[2][8] ), .IN2(n3605), .IN3(n3610), .IN4(n3801), 
        .Q(n522) );
  AO22X1 U2663 ( .IN1(\regfile[3][8] ), .IN2(n3597), .IN3(n3602), .IN4(n3801), 
        .Q(n521) );
  AO22X1 U2664 ( .IN1(\regfile[4][8] ), .IN2(n3589), .IN3(n3594), .IN4(n3801), 
        .Q(n520) );
  AO22X1 U2665 ( .IN1(\regfile[5][8] ), .IN2(n3581), .IN3(n3586), .IN4(n3801), 
        .Q(n519) );
  AO22X1 U2666 ( .IN1(\regfile[6][8] ), .IN2(n3573), .IN3(n3578), .IN4(n3801), 
        .Q(n518) );
  AO22X1 U2667 ( .IN1(\regfile[7][8] ), .IN2(n3565), .IN3(n3570), .IN4(n3801), 
        .Q(n517) );
  AO22X1 U2668 ( .IN1(\regfile[8][8] ), .IN2(n3557), .IN3(n3562), .IN4(n3801), 
        .Q(n516) );
  AO22X1 U2669 ( .IN1(\regfile[9][8] ), .IN2(n3549), .IN3(n3554), .IN4(n3801), 
        .Q(n515) );
  AO22X1 U2670 ( .IN1(\regfile[10][8] ), .IN2(n3541), .IN3(n3546), .IN4(n3801), 
        .Q(n514) );
  AO22X1 U2671 ( .IN1(\regfile[11][8] ), .IN2(n3533), .IN3(n3538), .IN4(n3801), 
        .Q(n513) );
  AO22X1 U2672 ( .IN1(\regfile[12][8] ), .IN2(n3525), .IN3(n3530), .IN4(n3801), 
        .Q(n512) );
  AO22X1 U2673 ( .IN1(\regfile[13][8] ), .IN2(n3517), .IN3(n3522), .IN4(n3801), 
        .Q(n511) );
  AO22X1 U2674 ( .IN1(\regfile[14][8] ), .IN2(n3509), .IN3(n3514), .IN4(n3801), 
        .Q(n510) );
  AO22X1 U2675 ( .IN1(\regfile[15][8] ), .IN2(n3501), .IN3(n3506), .IN4(n3801), 
        .Q(n509) );
  AO22X1 U2676 ( .IN1(\regfile[0][7] ), .IN2(n3621), .IN3(n3627), .IN4(n3802), 
        .Q(n508) );
  AO22X1 U2677 ( .IN1(\regfile[1][7] ), .IN2(n3613), .IN3(n3619), .IN4(n3802), 
        .Q(n507) );
  AO22X1 U2678 ( .IN1(\regfile[2][7] ), .IN2(n3605), .IN3(n3611), .IN4(n3802), 
        .Q(n506) );
  AO22X1 U2679 ( .IN1(\regfile[3][7] ), .IN2(n3597), .IN3(n3603), .IN4(n3802), 
        .Q(n505) );
  AO22X1 U2680 ( .IN1(\regfile[4][7] ), .IN2(n3589), .IN3(n3595), .IN4(n3802), 
        .Q(n504) );
  AO22X1 U2681 ( .IN1(\regfile[5][7] ), .IN2(n3581), .IN3(n3587), .IN4(n3802), 
        .Q(n503) );
  AO22X1 U2682 ( .IN1(\regfile[6][7] ), .IN2(n3573), .IN3(n3579), .IN4(n3802), 
        .Q(n502) );
  AO22X1 U2683 ( .IN1(\regfile[7][7] ), .IN2(n3565), .IN3(n3571), .IN4(n3802), 
        .Q(n501) );
  AO22X1 U2684 ( .IN1(\regfile[8][7] ), .IN2(n3557), .IN3(n3563), .IN4(n3802), 
        .Q(n500) );
  AO22X1 U2685 ( .IN1(\regfile[9][7] ), .IN2(n3549), .IN3(n3555), .IN4(n3802), 
        .Q(n499) );
  AO22X1 U2686 ( .IN1(\regfile[10][7] ), .IN2(n3541), .IN3(n3547), .IN4(n3802), 
        .Q(n498) );
  AO22X1 U2687 ( .IN1(\regfile[11][7] ), .IN2(n3533), .IN3(n3539), .IN4(n3802), 
        .Q(n497) );
  AO22X1 U2688 ( .IN1(\regfile[12][7] ), .IN2(n3525), .IN3(n3531), .IN4(n3802), 
        .Q(n496) );
  AO22X1 U2689 ( .IN1(\regfile[13][7] ), .IN2(n3517), .IN3(n3523), .IN4(n3802), 
        .Q(n495) );
  AO22X1 U2690 ( .IN1(\regfile[14][7] ), .IN2(n3509), .IN3(n3515), .IN4(n3802), 
        .Q(n494) );
  AO22X1 U2691 ( .IN1(\regfile[15][7] ), .IN2(n3501), .IN3(n3507), .IN4(n3802), 
        .Q(n493) );
  AO22X1 U2692 ( .IN1(\regfile[0][6] ), .IN2(n3621), .IN3(n3627), .IN4(n3803), 
        .Q(n492) );
  AO22X1 U2693 ( .IN1(\regfile[1][6] ), .IN2(n3613), .IN3(n3619), .IN4(n3803), 
        .Q(n491) );
  AO22X1 U2694 ( .IN1(\regfile[2][6] ), .IN2(n3605), .IN3(n3611), .IN4(n3803), 
        .Q(n490) );
  AO22X1 U2695 ( .IN1(\regfile[3][6] ), .IN2(n3597), .IN3(n3603), .IN4(n3803), 
        .Q(n489) );
  AO22X1 U2696 ( .IN1(\regfile[4][6] ), .IN2(n3589), .IN3(n3595), .IN4(n3803), 
        .Q(n488) );
  AO22X1 U2697 ( .IN1(\regfile[5][6] ), .IN2(n3581), .IN3(n3587), .IN4(n3803), 
        .Q(n487) );
  AO22X1 U2698 ( .IN1(\regfile[6][6] ), .IN2(n3573), .IN3(n3579), .IN4(n3803), 
        .Q(n486) );
  AO22X1 U2699 ( .IN1(\regfile[7][6] ), .IN2(n3565), .IN3(n3571), .IN4(n3803), 
        .Q(n485) );
  AO22X1 U2700 ( .IN1(\regfile[8][6] ), .IN2(n3557), .IN3(n3563), .IN4(n3803), 
        .Q(n484) );
  AO22X1 U2701 ( .IN1(\regfile[9][6] ), .IN2(n3549), .IN3(n3555), .IN4(n3803), 
        .Q(n483) );
  AO22X1 U2702 ( .IN1(\regfile[10][6] ), .IN2(n3541), .IN3(n3547), .IN4(n3803), 
        .Q(n482) );
  AO22X1 U2703 ( .IN1(\regfile[11][6] ), .IN2(n3533), .IN3(n3539), .IN4(n3803), 
        .Q(n481) );
  AO22X1 U2704 ( .IN1(\regfile[12][6] ), .IN2(n3525), .IN3(n3531), .IN4(n3803), 
        .Q(n480) );
  AO22X1 U2705 ( .IN1(\regfile[13][6] ), .IN2(n3517), .IN3(n3523), .IN4(n3803), 
        .Q(n479) );
  AO22X1 U2706 ( .IN1(\regfile[14][6] ), .IN2(n3509), .IN3(n3515), .IN4(n3803), 
        .Q(n478) );
  AO22X1 U2707 ( .IN1(\regfile[15][6] ), .IN2(n3501), .IN3(n3507), .IN4(n3803), 
        .Q(n477) );
  AO22X1 U2708 ( .IN1(\regfile[0][5] ), .IN2(n3621), .IN3(n3627), .IN4(n3804), 
        .Q(n476) );
  AO22X1 U2709 ( .IN1(\regfile[1][5] ), .IN2(n3613), .IN3(n3619), .IN4(n3804), 
        .Q(n475) );
  AO22X1 U2710 ( .IN1(\regfile[2][5] ), .IN2(n3605), .IN3(n3611), .IN4(n3804), 
        .Q(n474) );
  AO22X1 U2711 ( .IN1(\regfile[3][5] ), .IN2(n3597), .IN3(n3603), .IN4(n3804), 
        .Q(n473) );
  AO22X1 U2712 ( .IN1(\regfile[4][5] ), .IN2(n3589), .IN3(n3595), .IN4(n3804), 
        .Q(n472) );
  AO22X1 U2713 ( .IN1(\regfile[5][5] ), .IN2(n3581), .IN3(n3587), .IN4(n3804), 
        .Q(n471) );
  AO22X1 U2714 ( .IN1(\regfile[6][5] ), .IN2(n3573), .IN3(n3579), .IN4(n3804), 
        .Q(n470) );
  AO22X1 U2715 ( .IN1(\regfile[7][5] ), .IN2(n3565), .IN3(n3571), .IN4(n3804), 
        .Q(n469) );
  AO22X1 U2716 ( .IN1(\regfile[8][5] ), .IN2(n3557), .IN3(n3563), .IN4(n3804), 
        .Q(n468) );
  AO22X1 U2717 ( .IN1(\regfile[9][5] ), .IN2(n3549), .IN3(n3555), .IN4(n3804), 
        .Q(n467) );
  AO22X1 U2718 ( .IN1(\regfile[10][5] ), .IN2(n3541), .IN3(n3547), .IN4(n3804), 
        .Q(n466) );
  AO22X1 U2719 ( .IN1(\regfile[11][5] ), .IN2(n3533), .IN3(n3539), .IN4(n3804), 
        .Q(n465) );
  AO22X1 U2720 ( .IN1(\regfile[12][5] ), .IN2(n3525), .IN3(n3531), .IN4(n3804), 
        .Q(n464) );
  AO22X1 U2721 ( .IN1(\regfile[13][5] ), .IN2(n3517), .IN3(n3523), .IN4(n3804), 
        .Q(n463) );
  AO22X1 U2722 ( .IN1(\regfile[14][5] ), .IN2(n3509), .IN3(n3515), .IN4(n3804), 
        .Q(n462) );
  AO22X1 U2723 ( .IN1(\regfile[15][5] ), .IN2(n3501), .IN3(n3507), .IN4(n3804), 
        .Q(n461) );
  AO22X1 U2724 ( .IN1(\regfile[0][4] ), .IN2(n3621), .IN3(n3627), .IN4(n3805), 
        .Q(n460) );
  AO22X1 U2725 ( .IN1(\regfile[1][4] ), .IN2(n3613), .IN3(n3619), .IN4(n3805), 
        .Q(n459) );
  AO22X1 U2726 ( .IN1(\regfile[2][4] ), .IN2(n3605), .IN3(n3611), .IN4(n3805), 
        .Q(n458) );
  AO22X1 U2727 ( .IN1(\regfile[3][4] ), .IN2(n3597), .IN3(n3603), .IN4(n3805), 
        .Q(n457) );
  AO22X1 U2728 ( .IN1(\regfile[4][4] ), .IN2(n3589), .IN3(n3595), .IN4(n3805), 
        .Q(n456) );
  AO22X1 U2729 ( .IN1(\regfile[5][4] ), .IN2(n3581), .IN3(n3587), .IN4(n3805), 
        .Q(n455) );
  AO22X1 U2730 ( .IN1(\regfile[6][4] ), .IN2(n3573), .IN3(n3579), .IN4(n3805), 
        .Q(n454) );
  AO22X1 U2731 ( .IN1(\regfile[7][4] ), .IN2(n3565), .IN3(n3571), .IN4(n3805), 
        .Q(n453) );
  AO22X1 U2732 ( .IN1(\regfile[8][4] ), .IN2(n3557), .IN3(n3563), .IN4(n3805), 
        .Q(n452) );
  AO22X1 U2733 ( .IN1(\regfile[9][4] ), .IN2(n3549), .IN3(n3555), .IN4(n3805), 
        .Q(n451) );
  AO22X1 U2734 ( .IN1(\regfile[10][4] ), .IN2(n3541), .IN3(n3547), .IN4(n3805), 
        .Q(n450) );
  AO22X1 U2735 ( .IN1(\regfile[11][4] ), .IN2(n3533), .IN3(n3539), .IN4(n3805), 
        .Q(n449) );
  AO22X1 U2736 ( .IN1(\regfile[12][4] ), .IN2(n3525), .IN3(n3531), .IN4(n3805), 
        .Q(n448) );
  AO22X1 U2737 ( .IN1(\regfile[13][4] ), .IN2(n3517), .IN3(n3523), .IN4(n3805), 
        .Q(n447) );
  AO22X1 U2738 ( .IN1(\regfile[14][4] ), .IN2(n3509), .IN3(n3515), .IN4(n3805), 
        .Q(n446) );
  AO22X1 U2739 ( .IN1(\regfile[15][4] ), .IN2(n3501), .IN3(n3507), .IN4(n3805), 
        .Q(n445) );
  AO22X1 U2740 ( .IN1(\regfile[0][3] ), .IN2(n3620), .IN3(n3627), .IN4(n3806), 
        .Q(n444) );
  AO22X1 U2741 ( .IN1(\regfile[1][3] ), .IN2(n3612), .IN3(n3619), .IN4(n3806), 
        .Q(n443) );
  AO22X1 U2742 ( .IN1(\regfile[2][3] ), .IN2(n3604), .IN3(n3611), .IN4(n3806), 
        .Q(n442) );
  AO22X1 U2743 ( .IN1(\regfile[3][3] ), .IN2(n3596), .IN3(n3603), .IN4(n3806), 
        .Q(n441) );
  AO22X1 U2744 ( .IN1(\regfile[4][3] ), .IN2(n3588), .IN3(n3595), .IN4(n3806), 
        .Q(n440) );
  AO22X1 U2745 ( .IN1(\regfile[5][3] ), .IN2(n3580), .IN3(n3587), .IN4(n3806), 
        .Q(n439) );
  AO22X1 U2746 ( .IN1(\regfile[6][3] ), .IN2(n3572), .IN3(n3579), .IN4(n3806), 
        .Q(n438) );
  AO22X1 U2747 ( .IN1(\regfile[7][3] ), .IN2(n3564), .IN3(n3571), .IN4(n3806), 
        .Q(n437) );
  AO22X1 U2748 ( .IN1(\regfile[8][3] ), .IN2(n3556), .IN3(n3563), .IN4(n3806), 
        .Q(n436) );
  AO22X1 U2749 ( .IN1(\regfile[9][3] ), .IN2(n3548), .IN3(n3555), .IN4(n3806), 
        .Q(n435) );
  AO22X1 U2750 ( .IN1(\regfile[10][3] ), .IN2(n3540), .IN3(n3547), .IN4(n3806), 
        .Q(n434) );
  AO22X1 U2751 ( .IN1(\regfile[11][3] ), .IN2(n3532), .IN3(n3539), .IN4(n3806), 
        .Q(n433) );
  AO22X1 U2752 ( .IN1(\regfile[12][3] ), .IN2(n3524), .IN3(n3531), .IN4(n3806), 
        .Q(n432) );
  AO22X1 U2753 ( .IN1(\regfile[13][3] ), .IN2(n3516), .IN3(n3523), .IN4(n3806), 
        .Q(n431) );
  AO22X1 U2754 ( .IN1(\regfile[14][3] ), .IN2(n3508), .IN3(n3515), .IN4(n3806), 
        .Q(n430) );
  AO22X1 U2755 ( .IN1(\regfile[15][3] ), .IN2(n3500), .IN3(n3507), .IN4(n3806), 
        .Q(n429) );
  AO22X1 U2756 ( .IN1(\regfile[0][2] ), .IN2(n3620), .IN3(n3627), .IN4(n3807), 
        .Q(n428) );
  AO22X1 U2757 ( .IN1(\regfile[1][2] ), .IN2(n3612), .IN3(n3619), .IN4(n3807), 
        .Q(n427) );
  AO22X1 U2758 ( .IN1(\regfile[2][2] ), .IN2(n3604), .IN3(n3611), .IN4(n3807), 
        .Q(n426) );
  AO22X1 U2759 ( .IN1(\regfile[3][2] ), .IN2(n3596), .IN3(n3603), .IN4(n3807), 
        .Q(n425) );
  AO22X1 U2760 ( .IN1(\regfile[4][2] ), .IN2(n3588), .IN3(n3595), .IN4(n3807), 
        .Q(n424) );
  AO22X1 U2761 ( .IN1(\regfile[5][2] ), .IN2(n3580), .IN3(n3587), .IN4(n3807), 
        .Q(n423) );
  AO22X1 U2762 ( .IN1(\regfile[6][2] ), .IN2(n3572), .IN3(n3579), .IN4(n3807), 
        .Q(n422) );
  AO22X1 U2763 ( .IN1(\regfile[7][2] ), .IN2(n3564), .IN3(n3571), .IN4(n3807), 
        .Q(n421) );
  AO22X1 U2764 ( .IN1(\regfile[8][2] ), .IN2(n3556), .IN3(n3563), .IN4(n3807), 
        .Q(n420) );
  AO22X1 U2765 ( .IN1(\regfile[9][2] ), .IN2(n3548), .IN3(n3555), .IN4(n3807), 
        .Q(n419) );
  AO22X1 U2766 ( .IN1(\regfile[10][2] ), .IN2(n3540), .IN3(n3547), .IN4(n3807), 
        .Q(n418) );
  AO22X1 U2767 ( .IN1(\regfile[11][2] ), .IN2(n3532), .IN3(n3539), .IN4(n3807), 
        .Q(n417) );
  AO22X1 U2768 ( .IN1(\regfile[12][2] ), .IN2(n3524), .IN3(n3531), .IN4(n3807), 
        .Q(n416) );
  AO22X1 U2769 ( .IN1(\regfile[13][2] ), .IN2(n3516), .IN3(n3523), .IN4(n3807), 
        .Q(n415) );
  AO22X1 U2770 ( .IN1(\regfile[14][2] ), .IN2(n3508), .IN3(n3515), .IN4(n3807), 
        .Q(n414) );
  AO22X1 U2771 ( .IN1(\regfile[15][2] ), .IN2(n3500), .IN3(n3507), .IN4(n3807), 
        .Q(n413) );
  AO22X1 U2772 ( .IN1(\regfile[0][1] ), .IN2(n3620), .IN3(n3627), .IN4(n3808), 
        .Q(n412) );
  AO22X1 U2773 ( .IN1(\regfile[1][1] ), .IN2(n3612), .IN3(n3619), .IN4(n3808), 
        .Q(n411) );
  AO22X1 U2774 ( .IN1(\regfile[2][1] ), .IN2(n3604), .IN3(n3611), .IN4(n3808), 
        .Q(n410) );
  AO22X1 U2775 ( .IN1(\regfile[3][1] ), .IN2(n3596), .IN3(n3603), .IN4(n3808), 
        .Q(n409) );
  AO22X1 U2776 ( .IN1(\regfile[4][1] ), .IN2(n3588), .IN3(n3595), .IN4(n3808), 
        .Q(n408) );
  AO22X1 U2777 ( .IN1(\regfile[5][1] ), .IN2(n3580), .IN3(n3587), .IN4(n3808), 
        .Q(n407) );
  AO22X1 U2778 ( .IN1(\regfile[6][1] ), .IN2(n3572), .IN3(n3579), .IN4(n3808), 
        .Q(n406) );
  AO22X1 U2779 ( .IN1(\regfile[7][1] ), .IN2(n3564), .IN3(n3571), .IN4(n3808), 
        .Q(n405) );
  AO22X1 U2780 ( .IN1(\regfile[8][1] ), .IN2(n3556), .IN3(n3563), .IN4(n3808), 
        .Q(n404) );
  AO22X1 U2781 ( .IN1(\regfile[9][1] ), .IN2(n3548), .IN3(n3555), .IN4(n3808), 
        .Q(n403) );
  AO22X1 U2782 ( .IN1(\regfile[10][1] ), .IN2(n3540), .IN3(n3547), .IN4(n3808), 
        .Q(n402) );
  AO22X1 U2783 ( .IN1(\regfile[11][1] ), .IN2(n3532), .IN3(n3539), .IN4(n3808), 
        .Q(n401) );
  AO22X1 U2784 ( .IN1(\regfile[12][1] ), .IN2(n3524), .IN3(n3531), .IN4(n3808), 
        .Q(n400) );
  AO22X1 U2785 ( .IN1(\regfile[13][1] ), .IN2(n3516), .IN3(n3523), .IN4(n3808), 
        .Q(n399) );
  AO22X1 U2786 ( .IN1(\regfile[14][1] ), .IN2(n3508), .IN3(n3515), .IN4(n3808), 
        .Q(n398) );
  AO22X1 U2787 ( .IN1(\regfile[15][1] ), .IN2(n3500), .IN3(n3507), .IN4(n3808), 
        .Q(n397) );
  AO22X1 U2788 ( .IN1(\regfile[0][0] ), .IN2(n3620), .IN3(n3627), .IN4(n3809), 
        .Q(n396) );
  AO22X1 U2789 ( .IN1(\regfile[1][0] ), .IN2(n3612), .IN3(n3619), .IN4(n3809), 
        .Q(n395) );
  AO22X1 U2790 ( .IN1(\regfile[2][0] ), .IN2(n3604), .IN3(n3611), .IN4(n3809), 
        .Q(n394) );
  AO22X1 U2791 ( .IN1(\regfile[3][0] ), .IN2(n3596), .IN3(n3603), .IN4(n3809), 
        .Q(n393) );
  AO22X1 U2792 ( .IN1(\regfile[4][0] ), .IN2(n3588), .IN3(n3595), .IN4(n3809), 
        .Q(n392) );
  AO22X1 U2793 ( .IN1(\regfile[5][0] ), .IN2(n3580), .IN3(n3587), .IN4(n3809), 
        .Q(n391) );
  AO22X1 U2794 ( .IN1(\regfile[6][0] ), .IN2(n3572), .IN3(n3579), .IN4(n3809), 
        .Q(n390) );
  AO22X1 U2795 ( .IN1(\regfile[7][0] ), .IN2(n3564), .IN3(n3571), .IN4(n3809), 
        .Q(n389) );
  AO22X1 U2796 ( .IN1(\regfile[8][0] ), .IN2(n3556), .IN3(n3563), .IN4(n3809), 
        .Q(n388) );
  AO22X1 U2797 ( .IN1(\regfile[9][0] ), .IN2(n3548), .IN3(n3555), .IN4(n3809), 
        .Q(n387) );
  AO22X1 U2798 ( .IN1(\regfile[10][0] ), .IN2(n3540), .IN3(n3547), .IN4(n3809), 
        .Q(n386) );
  AO22X1 U2799 ( .IN1(\regfile[11][0] ), .IN2(n3532), .IN3(n3539), .IN4(n3809), 
        .Q(n385) );
  AO22X1 U2800 ( .IN1(\regfile[12][0] ), .IN2(n3524), .IN3(n3531), .IN4(n3809), 
        .Q(n384) );
  AO22X1 U2801 ( .IN1(\regfile[13][0] ), .IN2(n3516), .IN3(n3523), .IN4(n3809), 
        .Q(n383) );
  AND2X1 U2802 ( .IN1(n970), .IN2(n3224), .Q(n2843) );
  AO22X1 U2803 ( .IN1(\regfile[14][0] ), .IN2(n3508), .IN3(n3515), .IN4(n3809), 
        .Q(n382) );
  AND2X1 U2804 ( .IN1(n967), .IN2(n3225), .Q(n2845) );
  AO22X1 U2805 ( .IN1(\regfile[15][0] ), .IN2(n3500), .IN3(n3507), .IN4(n3809), 
        .Q(n381) );
  AND2X1 U2806 ( .IN1(n970), .IN2(n969), .Q(n2844) );
  AND2X1 U2807 ( .IN1(n967), .IN2(n968), .Q(n2846) );
  AND2X1 U2808 ( .IN1(n2847), .IN2(n2848), .Q(Zero) );
  NOR4X0 U2809 ( .IN1(n2849), .IN2(n2850), .IN3(n2851), .IN4(n2852), .QN(n2848) );
  NAND4X0 U2810 ( .IN1(n292), .IN2(n291), .IN3(n290), .IN4(n289), .QN(n2852)
         );
  NAND4X0 U2811 ( .IN1(n288), .IN2(n287), .IN3(n286), .IN4(n285), .QN(n2851)
         );
  NAND4X0 U2812 ( .IN1(n284), .IN2(n283), .IN3(n282), .IN4(n281), .QN(n2850)
         );
  NAND4X0 U2813 ( .IN1(n280), .IN2(n279), .IN3(n278), .IN4(n277), .QN(n2849)
         );
  NOR4X0 U2814 ( .IN1(n2853), .IN2(n2854), .IN3(n2855), .IN4(n2856), .QN(n2847) );
  NAND4X0 U2815 ( .IN1(n312), .IN2(n307), .IN3(n306), .IN4(n305), .QN(n2856)
         );
  NAND4X0 U2816 ( .IN1(n304), .IN2(n303), .IN3(n302), .IN4(n301), .QN(n2855)
         );
  NAND4X0 U2817 ( .IN1(n300), .IN2(n299), .IN3(n298), .IN4(n297), .QN(n2854)
         );
  NAND4X0 U2818 ( .IN1(n296), .IN2(n295), .IN3(n294), .IN4(n293), .QN(n2853)
         );
  OAI22X1 U2819 ( .IN1(n2857), .IN2(n2858), .IN3(n2859), .IN4(n2860), .QN(N325) );
  OA22X1 U2820 ( .IN1(n3810), .IN2(n2861), .IN3(n2862), .IN4(n3811), .Q(n2859)
         );
  AOI21X1 U2821 ( .IN1(n3810), .IN2(n344), .IN3(N257), .QN(n2862) );
  XNOR2X1 U2822 ( .IN1(N222), .IN2(N223), .Q(n2857) );
  AO22X1 U2823 ( .IN1(n3488), .IN2(N223), .IN3(N257), .IN4(n3486), .Q(N324) );
  AO221X1 U2824 ( .IN1(n3488), .IN2(N222), .IN3(n3499), .IN4(n3814), .IN5(
        n2864), .Q(N323) );
  AO222X1 U2825 ( .IN1(n2865), .IN2(n3810), .IN3(n2866), .IN4(n3483), .IN5(
        n3484), .IN6(N256), .Q(n2864) );
  AO21X1 U2826 ( .IN1(n3492), .IN2(n3814), .IN3(n3497), .Q(n2865) );
  AO221X1 U2827 ( .IN1(N221), .IN2(n3813), .IN3(n3499), .IN4(n3815), .IN5(
        n2868), .Q(N322) );
  AO222X1 U2828 ( .IN1(n2869), .IN2(IFID_B[30]), .IN3(n2870), .IN4(n379), 
        .IN5(N255), .IN6(n3484), .Q(n2868) );
  AO21X1 U2829 ( .IN1(n3492), .IN2(n3815), .IN3(n3497), .Q(n2869) );
  AO221X1 U2830 ( .IN1(N220), .IN2(n3813), .IN3(n3499), .IN4(n3816), .IN5(
        n2872), .Q(N321) );
  AO222X1 U2831 ( .IN1(n2873), .IN2(IFID_B[29]), .IN3(n2874), .IN4(n378), 
        .IN5(N254), .IN6(n3484), .Q(n2872) );
  AO21X1 U2832 ( .IN1(n3492), .IN2(n3816), .IN3(n3497), .Q(n2873) );
  AO221X1 U2833 ( .IN1(N219), .IN2(n3813), .IN3(n3499), .IN4(n3817), .IN5(
        n2875), .Q(N320) );
  AO222X1 U2834 ( .IN1(n2876), .IN2(IFID_B[28]), .IN3(n2877), .IN4(n377), 
        .IN5(N253), .IN6(n3484), .Q(n2875) );
  AO21X1 U2835 ( .IN1(n3492), .IN2(n3817), .IN3(n3497), .Q(n2876) );
  AO221X1 U2836 ( .IN1(N218), .IN2(n3813), .IN3(n3498), .IN4(n3818), .IN5(
        n2878), .Q(N319) );
  AO222X1 U2837 ( .IN1(n2879), .IN2(IFID_B[27]), .IN3(n2880), .IN4(n376), 
        .IN5(N252), .IN6(n3484), .Q(n2878) );
  AO21X1 U2838 ( .IN1(n3492), .IN2(n3818), .IN3(n3497), .Q(n2879) );
  AO221X1 U2839 ( .IN1(N217), .IN2(n3487), .IN3(n3498), .IN4(n3819), .IN5(
        n2881), .Q(N318) );
  AO222X1 U2840 ( .IN1(n2882), .IN2(IFID_B[26]), .IN3(n2883), .IN4(n375), 
        .IN5(N251), .IN6(n3484), .Q(n2881) );
  AO21X1 U2841 ( .IN1(n3492), .IN2(n3819), .IN3(n3497), .Q(n2882) );
  AO221X1 U2842 ( .IN1(N216), .IN2(n3488), .IN3(n3498), .IN4(n3820), .IN5(
        n2884), .Q(N317) );
  AO222X1 U2843 ( .IN1(n2885), .IN2(IFID_B[25]), .IN3(n2886), .IN4(n374), 
        .IN5(N250), .IN6(n3484), .Q(n2884) );
  AO21X1 U2844 ( .IN1(n3492), .IN2(n3820), .IN3(n3497), .Q(n2885) );
  AO221X1 U2845 ( .IN1(N215), .IN2(n3487), .IN3(n3498), .IN4(n3821), .IN5(
        n2887), .Q(N316) );
  AO222X1 U2846 ( .IN1(n2888), .IN2(IFID_B[24]), .IN3(n2889), .IN4(n373), 
        .IN5(N249), .IN6(n3485), .Q(n2887) );
  AO21X1 U2847 ( .IN1(n3492), .IN2(n3821), .IN3(n3496), .Q(n2888) );
  AO221X1 U2848 ( .IN1(N214), .IN2(n3488), .IN3(n3497), .IN4(n3822), .IN5(
        n2890), .Q(N315) );
  AO222X1 U2849 ( .IN1(n2891), .IN2(IFID_B[23]), .IN3(n2892), .IN4(n372), 
        .IN5(N248), .IN6(n3484), .Q(n2890) );
  AO21X1 U2850 ( .IN1(n3492), .IN2(n3822), .IN3(n3497), .Q(n2891) );
  AO221X1 U2851 ( .IN1(N213), .IN2(n3488), .IN3(n3498), .IN4(n3823), .IN5(
        n2893), .Q(N314) );
  AO222X1 U2852 ( .IN1(n2894), .IN2(IFID_B[22]), .IN3(n2895), .IN4(n371), 
        .IN5(N247), .IN6(n3484), .Q(n2893) );
  AO21X1 U2853 ( .IN1(n3492), .IN2(n3823), .IN3(n3496), .Q(n2894) );
  AO221X1 U2854 ( .IN1(N212), .IN2(n3488), .IN3(n3497), .IN4(n3824), .IN5(
        n2896), .Q(N313) );
  AO222X1 U2855 ( .IN1(n2897), .IN2(IFID_B[21]), .IN3(n2898), .IN4(n370), 
        .IN5(N246), .IN6(n3484), .Q(n2896) );
  AO21X1 U2856 ( .IN1(n3492), .IN2(n3824), .IN3(n3496), .Q(n2897) );
  AO221X1 U2857 ( .IN1(N211), .IN2(n3488), .IN3(n3497), .IN4(n3825), .IN5(
        n2899), .Q(N312) );
  AO222X1 U2858 ( .IN1(n2900), .IN2(IFID_B[20]), .IN3(n2901), .IN4(n369), 
        .IN5(N245), .IN6(n3484), .Q(n2899) );
  AO21X1 U2859 ( .IN1(n3492), .IN2(n3825), .IN3(n3496), .Q(n2900) );
  AO221X1 U2860 ( .IN1(N210), .IN2(n3488), .IN3(n3498), .IN4(n3826), .IN5(
        n2902), .Q(N311) );
  AO222X1 U2861 ( .IN1(n2903), .IN2(IFID_B[19]), .IN3(n2904), .IN4(n368), 
        .IN5(N244), .IN6(n3484), .Q(n2902) );
  AO21X1 U2862 ( .IN1(n3493), .IN2(n3826), .IN3(n3496), .Q(n2903) );
  AO221X1 U2863 ( .IN1(N209), .IN2(n3487), .IN3(n3497), .IN4(n3827), .IN5(
        n2905), .Q(N310) );
  AO222X1 U2864 ( .IN1(n2906), .IN2(IFID_B[18]), .IN3(n2907), .IN4(n367), 
        .IN5(N243), .IN6(n3484), .Q(n2905) );
  AO21X1 U2865 ( .IN1(n3493), .IN2(n3827), .IN3(n3496), .Q(n2906) );
  AO221X1 U2866 ( .IN1(N208), .IN2(n3487), .IN3(n3497), .IN4(n3828), .IN5(
        n2908), .Q(N309) );
  AO222X1 U2867 ( .IN1(n2909), .IN2(IFID_B[17]), .IN3(n2910), .IN4(n366), 
        .IN5(N242), .IN6(n3485), .Q(n2908) );
  AO21X1 U2868 ( .IN1(n3493), .IN2(n3828), .IN3(n3496), .Q(n2909) );
  AO221X1 U2869 ( .IN1(N207), .IN2(n3487), .IN3(n3498), .IN4(n3829), .IN5(
        n2911), .Q(N308) );
  AO222X1 U2870 ( .IN1(n2912), .IN2(IFID_B[16]), .IN3(n2913), .IN4(n365), 
        .IN5(N241), .IN6(n3485), .Q(n2911) );
  AO21X1 U2871 ( .IN1(n3493), .IN2(n3829), .IN3(n3496), .Q(n2912) );
  AO221X1 U2872 ( .IN1(N206), .IN2(n3487), .IN3(n3498), .IN4(n3830), .IN5(
        n2914), .Q(N307) );
  AO222X1 U2873 ( .IN1(n2915), .IN2(IFID_B[15]), .IN3(n2916), .IN4(n364), 
        .IN5(N240), .IN6(n3485), .Q(n2914) );
  AO21X1 U2874 ( .IN1(n3493), .IN2(n3830), .IN3(n3496), .Q(n2915) );
  AO221X1 U2875 ( .IN1(N205), .IN2(n3487), .IN3(n3498), .IN4(n3831), .IN5(
        n2917), .Q(N306) );
  AO222X1 U2876 ( .IN1(n2918), .IN2(IFID_B[14]), .IN3(n2919), .IN4(n363), 
        .IN5(N239), .IN6(n3485), .Q(n2917) );
  AO21X1 U2877 ( .IN1(n3493), .IN2(n3831), .IN3(n3496), .Q(n2918) );
  AO221X1 U2878 ( .IN1(N204), .IN2(n3487), .IN3(n3498), .IN4(n3832), .IN5(
        n2920), .Q(N305) );
  AO222X1 U2879 ( .IN1(n2921), .IN2(IFID_B[13]), .IN3(n2922), .IN4(n362), 
        .IN5(N238), .IN6(n3485), .Q(n2920) );
  AO21X1 U2880 ( .IN1(n3493), .IN2(n3832), .IN3(n3496), .Q(n2921) );
  AO221X1 U2881 ( .IN1(N203), .IN2(n3487), .IN3(n3498), .IN4(n3833), .IN5(
        n2923), .Q(N304) );
  AO222X1 U2882 ( .IN1(n2924), .IN2(IFID_B[12]), .IN3(n2925), .IN4(n361), 
        .IN5(N237), .IN6(n3485), .Q(n2923) );
  AO21X1 U2883 ( .IN1(n3493), .IN2(n3833), .IN3(n3495), .Q(n2924) );
  AO221X1 U2884 ( .IN1(N202), .IN2(n3487), .IN3(n3498), .IN4(n3834), .IN5(
        n2926), .Q(N303) );
  AO222X1 U2885 ( .IN1(n2927), .IN2(IFID_B[11]), .IN3(n2928), .IN4(n360), 
        .IN5(N236), .IN6(n3485), .Q(n2926) );
  AO21X1 U2886 ( .IN1(n3493), .IN2(n3834), .IN3(n3495), .Q(n2927) );
  AO221X1 U2887 ( .IN1(N201), .IN2(n3487), .IN3(n3499), .IN4(n3835), .IN5(
        n2929), .Q(N302) );
  AO222X1 U2888 ( .IN1(n2930), .IN2(IFID_B[10]), .IN3(n2931), .IN4(n359), 
        .IN5(N235), .IN6(n3485), .Q(n2929) );
  AO21X1 U2889 ( .IN1(n3493), .IN2(n3835), .IN3(n3495), .Q(n2930) );
  AO221X1 U2890 ( .IN1(N200), .IN2(n3487), .IN3(n3498), .IN4(n3836), .IN5(
        n2932), .Q(N301) );
  AO222X1 U2891 ( .IN1(n2933), .IN2(IFID_B[9]), .IN3(n2934), .IN4(n358), .IN5(
        N234), .IN6(n3485), .Q(n2932) );
  AO21X1 U2892 ( .IN1(n3493), .IN2(n3836), .IN3(n3495), .Q(n2933) );
  AO221X1 U2893 ( .IN1(N199), .IN2(n3487), .IN3(n3498), .IN4(n3837), .IN5(
        n2935), .Q(N300) );
  AO222X1 U2894 ( .IN1(n2936), .IN2(IFID_B[8]), .IN3(n2937), .IN4(n357), .IN5(
        N233), .IN6(n3485), .Q(n2935) );
  AO21X1 U2895 ( .IN1(n3493), .IN2(n3837), .IN3(n3495), .Q(n2936) );
  AO221X1 U2896 ( .IN1(N198), .IN2(n3487), .IN3(n3499), .IN4(n3838), .IN5(
        n2938), .Q(N299) );
  AO222X1 U2897 ( .IN1(n2939), .IN2(IFID_B[7]), .IN3(n2940), .IN4(n356), .IN5(
        N232), .IN6(n3485), .Q(n2938) );
  AO21X1 U2898 ( .IN1(n3494), .IN2(n3838), .IN3(n3495), .Q(n2939) );
  AO221X1 U2899 ( .IN1(N197), .IN2(n3487), .IN3(n3499), .IN4(n3839), .IN5(
        n2941), .Q(N298) );
  AO222X1 U2900 ( .IN1(n2942), .IN2(IFID_B[6]), .IN3(n2943), .IN4(n355), .IN5(
        N231), .IN6(n3485), .Q(n2941) );
  AO21X1 U2901 ( .IN1(n3494), .IN2(n3839), .IN3(n3495), .Q(n2942) );
  AO221X1 U2902 ( .IN1(N196), .IN2(n3488), .IN3(n3499), .IN4(n3840), .IN5(
        n2944), .Q(N297) );
  AO222X1 U2903 ( .IN1(n2945), .IN2(IFID_B[5]), .IN3(n2946), .IN4(n354), .IN5(
        N230), .IN6(n3486), .Q(n2944) );
  AO21X1 U2904 ( .IN1(n3494), .IN2(n3840), .IN3(n3495), .Q(n2945) );
  AO221X1 U2905 ( .IN1(N195), .IN2(n3488), .IN3(n3499), .IN4(n3841), .IN5(
        n2947), .Q(N296) );
  AO222X1 U2906 ( .IN1(n2948), .IN2(IFID_B[4]), .IN3(n2949), .IN4(n353), .IN5(
        N229), .IN6(n3486), .Q(n2947) );
  AO21X1 U2907 ( .IN1(n3494), .IN2(n3841), .IN3(n3495), .Q(n2948) );
  AO221X1 U2908 ( .IN1(N194), .IN2(n3488), .IN3(n3499), .IN4(n3842), .IN5(
        n2950), .Q(N295) );
  AO222X1 U2909 ( .IN1(n2951), .IN2(IFID_B[3]), .IN3(n2952), .IN4(n352), .IN5(
        N228), .IN6(n3486), .Q(n2950) );
  AO21X1 U2910 ( .IN1(n3494), .IN2(n3842), .IN3(n3495), .Q(n2951) );
  AO221X1 U2911 ( .IN1(N193), .IN2(n3488), .IN3(n3499), .IN4(n3843), .IN5(
        n2953), .Q(N294) );
  AO222X1 U2912 ( .IN1(n2954), .IN2(IFID_B[2]), .IN3(n2955), .IN4(n351), .IN5(
        N227), .IN6(n3486), .Q(n2953) );
  AO21X1 U2913 ( .IN1(n3494), .IN2(n3843), .IN3(n3495), .Q(n2954) );
  AO221X1 U2914 ( .IN1(N192), .IN2(n3813), .IN3(n3499), .IN4(n3844), .IN5(
        n2956), .Q(N293) );
  AO222X1 U2915 ( .IN1(n2957), .IN2(IFID_B[1]), .IN3(n2958), .IN4(n350), .IN5(
        N226), .IN6(n3486), .Q(n2956) );
  AO21X1 U2916 ( .IN1(n3494), .IN2(n3844), .IN3(n3495), .Q(n2957) );
  NAND4X0 U2917 ( .IN1(n2959), .IN2(n2960), .IN3(n2961), .IN4(n2962), .QN(N292) );
  AOI222X1 U2918 ( .IN1(n3499), .IN2(n3845), .IN3(N225), .IN4(n3486), .IN5(
        N191), .IN6(n3813), .QN(n2962) );
  NOR3X0 U2919 ( .IN1(n971), .IN2(n972), .IN3(n2966), .QN(n2963) );
  AO21X1 U2920 ( .IN1(n3494), .IN2(n3845), .IN3(n3496), .Q(n2964) );
  AND2X1 U2921 ( .IN1(n3494), .IN2(n971), .Q(n2863) );
  NOR3X0 U2922 ( .IN1(n972), .IN2(n973), .IN3(n966), .QN(n2867) );
  NAND4X0 U2923 ( .IN1(N259), .IN2(n971), .IN3(n2965), .IN4(n973), .QN(n2960)
         );
  NAND3X0 U2924 ( .IN1(n313), .IN2(n3483), .IN3(n349), .QN(n2959) );
  pipealu_DW_cmp_0 lt_85 ( .A(IFID_A), .B(IFID_B), .TC(1'b0), .GE_LT(1'b1), 
        .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N259) );
  pipealu_DW01_sub_0 sub_78 ( .A({1'b0, IFID_A}), .B({1'b0, IFID_B}), .CI(1'b0), .DIFF({N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, 
        N234, N233, N232, N231, N230, N229, N228, N227, N226, N225}) );
  pipealu_DW01_add_0 add_73 ( .A({1'b0, IFID_A}), .B({1'b0, IFID_B}), .CI(1'b0), .SUM({N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, 
        N199, N198, N197, N196, N195, N194, N193, N192, N191}) );
  INVX0 U2926 ( .INP(rst), .ZN(n3769) );
  NBUFFX2 U2927 ( .INP(n3813), .Z(n3488) );
  INVX0 U2928 ( .INP(n3500), .ZN(n3506) );
  INVX0 U2929 ( .INP(n3508), .ZN(n3514) );
  INVX0 U2930 ( .INP(n3516), .ZN(n3522) );
  INVX0 U2931 ( .INP(n3524), .ZN(n3530) );
  INVX0 U2932 ( .INP(n3532), .ZN(n3538) );
  INVX0 U2933 ( .INP(n3540), .ZN(n3546) );
  INVX0 U2934 ( .INP(n3548), .ZN(n3554) );
  INVX0 U2935 ( .INP(n3556), .ZN(n3562) );
  INVX0 U2936 ( .INP(n3564), .ZN(n3570) );
  INVX0 U2937 ( .INP(n3572), .ZN(n3578) );
  INVX0 U2938 ( .INP(n3580), .ZN(n3586) );
  INVX0 U2939 ( .INP(n3588), .ZN(n3594) );
  INVX0 U2940 ( .INP(n3596), .ZN(n3602) );
  INVX0 U2941 ( .INP(n3604), .ZN(n3610) );
  INVX0 U2942 ( .INP(n3612), .ZN(n3618) );
  INVX0 U2943 ( .INP(n3620), .ZN(n3626) );
  INVX0 U2944 ( .INP(n3500), .ZN(n3505) );
  INVX0 U2945 ( .INP(n3508), .ZN(n3513) );
  INVX0 U2946 ( .INP(n3516), .ZN(n3521) );
  INVX0 U2947 ( .INP(n3524), .ZN(n3529) );
  INVX0 U2948 ( .INP(n3532), .ZN(n3537) );
  INVX0 U2949 ( .INP(n3540), .ZN(n3545) );
  INVX0 U2950 ( .INP(n3548), .ZN(n3553) );
  INVX0 U2951 ( .INP(n3556), .ZN(n3561) );
  INVX0 U2952 ( .INP(n3564), .ZN(n3569) );
  INVX0 U2953 ( .INP(n3572), .ZN(n3577) );
  INVX0 U2954 ( .INP(n3580), .ZN(n3585) );
  INVX0 U2955 ( .INP(n3588), .ZN(n3593) );
  INVX0 U2956 ( .INP(n3596), .ZN(n3601) );
  INVX0 U2957 ( .INP(n3604), .ZN(n3609) );
  INVX0 U2958 ( .INP(n3612), .ZN(n3617) );
  INVX0 U2959 ( .INP(n3620), .ZN(n3625) );
  NBUFFX2 U2960 ( .INP(n2219), .Z(n3687) );
  NBUFFX2 U2961 ( .INP(n2531), .Z(n3639) );
  NBUFFX2 U2962 ( .INP(n2838), .Z(n3500) );
  NBUFFX2 U2963 ( .INP(n2837), .Z(n3508) );
  NBUFFX2 U2964 ( .INP(n2836), .Z(n3516) );
  NBUFFX2 U2965 ( .INP(n2835), .Z(n3524) );
  NBUFFX2 U2966 ( .INP(n2834), .Z(n3532) );
  NBUFFX2 U2967 ( .INP(n2833), .Z(n3540) );
  NBUFFX2 U2968 ( .INP(n2832), .Z(n3548) );
  NBUFFX2 U2969 ( .INP(n2831), .Z(n3556) );
  NBUFFX2 U2970 ( .INP(n2830), .Z(n3564) );
  NBUFFX2 U2971 ( .INP(n2829), .Z(n3572) );
  NBUFFX2 U2972 ( .INP(n2828), .Z(n3580) );
  NBUFFX2 U2973 ( .INP(n2827), .Z(n3588) );
  NBUFFX2 U2974 ( .INP(n2826), .Z(n3596) );
  NBUFFX2 U2975 ( .INP(n2825), .Z(n3604) );
  NBUFFX2 U2976 ( .INP(n2824), .Z(n3612) );
  NBUFFX2 U2977 ( .INP(n2823), .Z(n3620) );
  NBUFFX2 U2978 ( .INP(n3812), .Z(n3486) );
  NBUFFX2 U2979 ( .INP(n2826), .Z(n3597) );
  NBUFFX2 U2980 ( .INP(n2825), .Z(n3605) );
  NBUFFX2 U2981 ( .INP(n2824), .Z(n3613) );
  NBUFFX2 U2982 ( .INP(n2823), .Z(n3621) );
  NBUFFX2 U2983 ( .INP(n2826), .Z(n3598) );
  NBUFFX2 U2984 ( .INP(n2825), .Z(n3606) );
  NBUFFX2 U2985 ( .INP(n2824), .Z(n3614) );
  NBUFFX2 U2986 ( .INP(n2823), .Z(n3622) );
  NBUFFX2 U2987 ( .INP(n2826), .Z(n3599) );
  NBUFFX2 U2988 ( .INP(n2825), .Z(n3607) );
  NBUFFX2 U2989 ( .INP(n2824), .Z(n3615) );
  NBUFFX2 U2990 ( .INP(n2823), .Z(n3623) );
  NBUFFX2 U2991 ( .INP(n2826), .Z(n3600) );
  NBUFFX2 U2992 ( .INP(n2825), .Z(n3608) );
  NBUFFX2 U2993 ( .INP(n2824), .Z(n3616) );
  NBUFFX2 U2994 ( .INP(n2823), .Z(n3624) );
  NBUFFX2 U2995 ( .INP(n2838), .Z(n3501) );
  NBUFFX2 U2996 ( .INP(n2837), .Z(n3509) );
  NBUFFX2 U2997 ( .INP(n2836), .Z(n3517) );
  NBUFFX2 U2998 ( .INP(n2835), .Z(n3525) );
  NBUFFX2 U2999 ( .INP(n2834), .Z(n3533) );
  NBUFFX2 U3000 ( .INP(n2833), .Z(n3541) );
  NBUFFX2 U3001 ( .INP(n2832), .Z(n3549) );
  NBUFFX2 U3002 ( .INP(n2831), .Z(n3557) );
  NBUFFX2 U3003 ( .INP(n2830), .Z(n3565) );
  NBUFFX2 U3004 ( .INP(n2829), .Z(n3573) );
  NBUFFX2 U3005 ( .INP(n2828), .Z(n3581) );
  NBUFFX2 U3006 ( .INP(n2827), .Z(n3589) );
  NBUFFX2 U3007 ( .INP(n2838), .Z(n3502) );
  NBUFFX2 U3008 ( .INP(n2837), .Z(n3510) );
  NBUFFX2 U3009 ( .INP(n2836), .Z(n3518) );
  NBUFFX2 U3010 ( .INP(n2835), .Z(n3526) );
  NBUFFX2 U3011 ( .INP(n2834), .Z(n3534) );
  NBUFFX2 U3012 ( .INP(n2833), .Z(n3542) );
  NBUFFX2 U3013 ( .INP(n2832), .Z(n3550) );
  NBUFFX2 U3014 ( .INP(n2831), .Z(n3558) );
  NBUFFX2 U3015 ( .INP(n2830), .Z(n3566) );
  NBUFFX2 U3016 ( .INP(n2829), .Z(n3574) );
  NBUFFX2 U3017 ( .INP(n2828), .Z(n3582) );
  NBUFFX2 U3018 ( .INP(n2827), .Z(n3590) );
  NBUFFX2 U3019 ( .INP(n2838), .Z(n3503) );
  NBUFFX2 U3020 ( .INP(n2837), .Z(n3511) );
  NBUFFX2 U3021 ( .INP(n2836), .Z(n3519) );
  NBUFFX2 U3022 ( .INP(n2835), .Z(n3527) );
  NBUFFX2 U3023 ( .INP(n2834), .Z(n3535) );
  NBUFFX2 U3024 ( .INP(n2833), .Z(n3543) );
  NBUFFX2 U3025 ( .INP(n2832), .Z(n3551) );
  NBUFFX2 U3026 ( .INP(n2831), .Z(n3559) );
  NBUFFX2 U3027 ( .INP(n2830), .Z(n3567) );
  NBUFFX2 U3028 ( .INP(n2829), .Z(n3575) );
  NBUFFX2 U3029 ( .INP(n2828), .Z(n3583) );
  NBUFFX2 U3030 ( .INP(n2827), .Z(n3591) );
  NBUFFX2 U3031 ( .INP(n2838), .Z(n3504) );
  NBUFFX2 U3032 ( .INP(n2837), .Z(n3512) );
  NBUFFX2 U3033 ( .INP(n2836), .Z(n3520) );
  NBUFFX2 U3034 ( .INP(n2835), .Z(n3528) );
  NBUFFX2 U3035 ( .INP(n2834), .Z(n3536) );
  NBUFFX2 U3036 ( .INP(n2833), .Z(n3544) );
  NBUFFX2 U3037 ( .INP(n2832), .Z(n3552) );
  NBUFFX2 U3038 ( .INP(n2831), .Z(n3560) );
  NBUFFX2 U3039 ( .INP(n2830), .Z(n3568) );
  NBUFFX2 U3040 ( .INP(n2829), .Z(n3576) );
  NBUFFX2 U3041 ( .INP(n2828), .Z(n3584) );
  NBUFFX2 U3042 ( .INP(n2827), .Z(n3592) );
  INVX0 U3043 ( .INP(n2858), .ZN(n3813) );
  NBUFFX2 U3044 ( .INP(n2519), .Z(n3669) );
  NBUFFX2 U3045 ( .INP(n2524), .Z(n3657) );
  NBUFFX2 U3046 ( .INP(n2529), .Z(n3645) );
  NBUFFX2 U3047 ( .INP(n2534), .Z(n3633) );
  NBUFFX2 U3048 ( .INP(n2207), .Z(n3717) );
  NBUFFX2 U3049 ( .INP(n2212), .Z(n3705) );
  NBUFFX2 U3050 ( .INP(n2217), .Z(n3693) );
  NBUFFX2 U3051 ( .INP(n2222), .Z(n3681) );
  NBUFFX2 U3052 ( .INP(n2520), .Z(n3666) );
  NBUFFX2 U3053 ( .INP(n2525), .Z(n3654) );
  NBUFFX2 U3054 ( .INP(n2530), .Z(n3642) );
  NBUFFX2 U3055 ( .INP(n2535), .Z(n3630) );
  NBUFFX2 U3056 ( .INP(n2208), .Z(n3714) );
  NBUFFX2 U3057 ( .INP(n2213), .Z(n3702) );
  NBUFFX2 U3058 ( .INP(n2218), .Z(n3690) );
  NBUFFX2 U3059 ( .INP(n2223), .Z(n3678) );
  NBUFFX2 U3060 ( .INP(n2204), .Z(n3723) );
  NBUFFX2 U3061 ( .INP(n2209), .Z(n3711) );
  NBUFFX2 U3062 ( .INP(n2214), .Z(n3699) );
  NBUFFX2 U3063 ( .INP(n2517), .Z(n3672) );
  NBUFFX2 U3064 ( .INP(n2522), .Z(n3660) );
  NBUFFX2 U3065 ( .INP(n2527), .Z(n3648) );
  NBUFFX2 U3066 ( .INP(n2532), .Z(n3636) );
  NBUFFX2 U3067 ( .INP(n2205), .Z(n3720) );
  NBUFFX2 U3068 ( .INP(n2210), .Z(n3708) );
  NBUFFX2 U3069 ( .INP(n2215), .Z(n3696) );
  NBUFFX2 U3070 ( .INP(n2220), .Z(n3684) );
  NBUFFX2 U3071 ( .INP(n2521), .Z(n3663) );
  NBUFFX2 U3072 ( .INP(n2526), .Z(n3651) );
  NBUFFX2 U3073 ( .INP(n2516), .Z(n3675) );
  NAND2X1 U3074 ( .IN1(n2822), .IN2(n2816), .QN(n2531) );
  NAND2X1 U3075 ( .IN1(n2510), .IN2(n2504), .QN(n2219) );
  NOR2X0 U3076 ( .IN1(n3810), .IN2(n3814), .QN(n2866) );
  INVX0 U3077 ( .INP(N256), .ZN(n3811) );
  NAND2X1 U3078 ( .IN1(n3811), .IN2(n3814), .QN(n2861) );
  INVX0 U3079 ( .INP(n3483), .ZN(n3489) );
  INVX0 U3080 ( .INP(n3483), .ZN(n3490) );
  NAND2X1 U3081 ( .IN1(n2963), .IN2(n3223), .QN(n2858) );
  NAND2X1 U3082 ( .IN1(n2846), .IN2(n2844), .QN(n2838) );
  NAND2X1 U3083 ( .IN1(n2845), .IN2(n2844), .QN(n2837) );
  NAND2X1 U3084 ( .IN1(n2846), .IN2(n2843), .QN(n2836) );
  NAND2X1 U3085 ( .IN1(n2845), .IN2(n2843), .QN(n2835) );
  NAND2X1 U3086 ( .IN1(n2846), .IN2(n2842), .QN(n2834) );
  NAND2X1 U3087 ( .IN1(n2845), .IN2(n2842), .QN(n2833) );
  NAND2X1 U3088 ( .IN1(n2844), .IN2(n2841), .QN(n2830) );
  NAND2X1 U3089 ( .IN1(n2844), .IN2(n2839), .QN(n2829) );
  NAND2X1 U3090 ( .IN1(n2843), .IN2(n2841), .QN(n2828) );
  NAND2X1 U3091 ( .IN1(n2843), .IN2(n2839), .QN(n2827) );
  NAND2X1 U3092 ( .IN1(n2842), .IN2(n2841), .QN(n2826) );
  NAND2X1 U3093 ( .IN1(n2842), .IN2(n2839), .QN(n2825) );
  INVX0 U3094 ( .INP(n2860), .ZN(n3812) );
  NAND2X1 U3095 ( .IN1(n2846), .IN2(n2840), .QN(n2832) );
  NAND2X1 U3096 ( .IN1(n2845), .IN2(n2840), .QN(n2831) );
  NAND2X1 U3097 ( .IN1(n2841), .IN2(n2840), .QN(n2824) );
  NAND2X1 U3098 ( .IN1(n2839), .IN2(n2840), .QN(n2823) );
  NOR2X0 U3099 ( .IN1(n3848), .IN2(n3849), .QN(n2816) );
  NOR2X0 U3100 ( .IN1(n3852), .IN2(n3853), .QN(n2504) );
  NOR2X0 U3101 ( .IN1(n3846), .IN2(n3847), .QN(n2822) );
  NOR2X0 U3102 ( .IN1(n3850), .IN2(n3851), .QN(n2510) );
  NAND2X1 U3103 ( .IN1(n2818), .IN2(n2816), .QN(n2521) );
  NAND2X1 U3104 ( .IN1(n2820), .IN2(n2816), .QN(n2526) );
  NAND2X1 U3105 ( .IN1(n2506), .IN2(n2504), .QN(n2209) );
  NAND2X1 U3106 ( .IN1(n2508), .IN2(n2504), .QN(n2214) );
  NAND2X1 U3107 ( .IN1(n2812), .IN2(n2813), .QN(n2520) );
  NAND2X1 U3108 ( .IN1(n2818), .IN2(n2812), .QN(n2525) );
  NAND2X1 U3109 ( .IN1(n2820), .IN2(n2812), .QN(n2530) );
  NAND2X1 U3110 ( .IN1(n2822), .IN2(n2812), .QN(n2535) );
  NAND2X1 U3111 ( .IN1(n2500), .IN2(n2501), .QN(n2208) );
  NAND2X1 U3112 ( .IN1(n2506), .IN2(n2500), .QN(n2213) );
  NAND2X1 U3113 ( .IN1(n2508), .IN2(n2500), .QN(n2218) );
  NAND2X1 U3114 ( .IN1(n2510), .IN2(n2500), .QN(n2223) );
  NAND2X1 U3115 ( .IN1(n2815), .IN2(n2813), .QN(n2517) );
  NAND2X1 U3116 ( .IN1(n2816), .IN2(n2813), .QN(n2516) );
  NAND2X1 U3117 ( .IN1(n2818), .IN2(n2815), .QN(n2522) );
  NAND2X1 U3118 ( .IN1(n2820), .IN2(n2815), .QN(n2527) );
  NAND2X1 U3119 ( .IN1(n2822), .IN2(n2815), .QN(n2532) );
  NAND2X1 U3120 ( .IN1(n2504), .IN2(n2501), .QN(n2204) );
  NAND2X1 U3121 ( .IN1(n2503), .IN2(n2501), .QN(n2205) );
  NAND2X1 U3122 ( .IN1(n2506), .IN2(n2503), .QN(n2210) );
  NAND2X1 U3123 ( .IN1(n2508), .IN2(n2503), .QN(n2215) );
  NAND2X1 U3124 ( .IN1(n2510), .IN2(n2503), .QN(n2220) );
  NAND2X1 U3125 ( .IN1(n2813), .IN2(n2814), .QN(n2519) );
  NAND2X1 U3126 ( .IN1(n2818), .IN2(n2814), .QN(n2524) );
  NAND2X1 U3127 ( .IN1(n2820), .IN2(n2814), .QN(n2529) );
  NAND2X1 U3128 ( .IN1(n2822), .IN2(n2814), .QN(n2534) );
  NAND2X1 U3129 ( .IN1(n2501), .IN2(n2502), .QN(n2207) );
  NAND2X1 U3130 ( .IN1(n2506), .IN2(n2502), .QN(n2212) );
  NAND2X1 U3131 ( .IN1(n2508), .IN2(n2502), .QN(n2217) );
  NAND2X1 U3132 ( .IN1(n2510), .IN2(n2502), .QN(n2222) );
  INVX0 U3133 ( .INP(n3769), .ZN(n3765) );
  INVX0 U3134 ( .INP(n3769), .ZN(n3766) );
  INVX0 U3135 ( .INP(n3769), .ZN(n3767) );
  INVX0 U3136 ( .INP(n3769), .ZN(n3768) );
  NOR2X0 U3137 ( .IN1(n3491), .IN2(n3818), .QN(n2880) );
  NOR2X0 U3138 ( .IN1(n3491), .IN2(n3817), .QN(n2877) );
  NOR2X0 U3139 ( .IN1(n3491), .IN2(n3816), .QN(n2874) );
  NOR2X0 U3140 ( .IN1(n3491), .IN2(n3815), .QN(n2870) );
  NOR2X0 U3141 ( .IN1(n3490), .IN2(n3828), .QN(n2910) );
  NOR2X0 U3142 ( .IN1(n3490), .IN2(n3826), .QN(n2904) );
  NOR2X0 U3143 ( .IN1(n3490), .IN2(n3824), .QN(n2898) );
  NOR2X0 U3144 ( .IN1(n3490), .IN2(n3822), .QN(n2892) );
  NOR2X0 U3145 ( .IN1(n3490), .IN2(n3821), .QN(n2889) );
  NOR2X0 U3146 ( .IN1(n3490), .IN2(n3827), .QN(n2907) );
  NOR2X0 U3147 ( .IN1(n3490), .IN2(n3823), .QN(n2895) );
  NOR2X0 U3148 ( .IN1(n3491), .IN2(n3820), .QN(n2886) );
  NOR2X0 U3149 ( .IN1(n3491), .IN2(n3819), .QN(n2883) );
  NOR2X0 U3150 ( .IN1(n3490), .IN2(n3825), .QN(n2901) );
  NOR2X0 U3151 ( .IN1(n3489), .IN2(n3838), .QN(n2940) );
  NOR2X0 U3152 ( .IN1(n3489), .IN2(n3837), .QN(n2937) );
  NOR2X0 U3153 ( .IN1(n3489), .IN2(n3834), .QN(n2928) );
  NOR2X0 U3154 ( .IN1(n3489), .IN2(n3833), .QN(n2925) );
  NOR2X0 U3155 ( .IN1(n3490), .IN2(n3830), .QN(n2916) );
  NOR2X0 U3156 ( .IN1(n3489), .IN2(n3839), .QN(n2943) );
  NOR2X0 U3157 ( .IN1(n3489), .IN2(n3836), .QN(n2934) );
  NOR2X0 U3158 ( .IN1(n3489), .IN2(n3835), .QN(n2931) );
  NOR2X0 U3159 ( .IN1(n3490), .IN2(n3832), .QN(n2922) );
  NOR2X0 U3160 ( .IN1(n3490), .IN2(n3831), .QN(n2919) );
  NOR2X0 U3161 ( .IN1(n3490), .IN2(n3829), .QN(n2913) );
  AND4X1 U3162 ( .IN1(n966), .IN2(n972), .IN3(n3482), .IN4(n2966), .Q(n3483)
         );
  NOR2X0 U3163 ( .IN1(n970), .IN2(n969), .QN(n2840) );
  NOR2X0 U3164 ( .IN1(n968), .IN2(n967), .QN(n2839) );
  NOR2X0 U3165 ( .IN1(n3225), .IN2(n967), .QN(n2841) );
  NOR2X0 U3166 ( .IN1(n3224), .IN2(n970), .QN(n2842) );
  INVX0 U3167 ( .INP(n344), .ZN(n3814) );
  INVX0 U3168 ( .INP(n279), .ZN(n3807) );
  INVX0 U3169 ( .INP(n283), .ZN(n3803) );
  INVX0 U3170 ( .INP(n287), .ZN(n3799) );
  INVX0 U3171 ( .INP(n291), .ZN(n3795) );
  INVX0 U3172 ( .INP(n295), .ZN(n3791) );
  INVX0 U3173 ( .INP(n299), .ZN(n3787) );
  INVX0 U3174 ( .INP(n303), .ZN(n3783) );
  INVX0 U3175 ( .INP(n307), .ZN(n3779) );
  INVX0 U3176 ( .INP(n280), .ZN(n3806) );
  INVX0 U3177 ( .INP(n284), .ZN(n3802) );
  INVX0 U3178 ( .INP(n288), .ZN(n3798) );
  INVX0 U3179 ( .INP(n292), .ZN(n3794) );
  INVX0 U3180 ( .INP(n296), .ZN(n3790) );
  INVX0 U3181 ( .INP(n300), .ZN(n3786) );
  INVX0 U3182 ( .INP(n304), .ZN(n3782) );
  INVX0 U3183 ( .INP(n312), .ZN(n3778) );
  INVX0 U3184 ( .INP(n278), .ZN(n3808) );
  INVX0 U3185 ( .INP(n282), .ZN(n3804) );
  INVX0 U3186 ( .INP(n286), .ZN(n3800) );
  INVX0 U3187 ( .INP(n290), .ZN(n3796) );
  INVX0 U3188 ( .INP(n294), .ZN(n3792) );
  INVX0 U3189 ( .INP(n298), .ZN(n3788) );
  INVX0 U3190 ( .INP(n302), .ZN(n3784) );
  INVX0 U3191 ( .INP(n306), .ZN(n3780) );
  INVX0 U3192 ( .INP(n277), .ZN(n3809) );
  INVX0 U3193 ( .INP(n281), .ZN(n3805) );
  INVX0 U3194 ( .INP(n285), .ZN(n3801) );
  INVX0 U3195 ( .INP(n289), .ZN(n3797) );
  INVX0 U3196 ( .INP(n293), .ZN(n3793) );
  INVX0 U3197 ( .INP(n297), .ZN(n3789) );
  INVX0 U3198 ( .INP(n301), .ZN(n3785) );
  INVX0 U3199 ( .INP(n305), .ZN(n3781) );
  NAND2X1 U3200 ( .IN1(n2964), .IN2(IFID_B[0]), .QN(n2961) );
  INVX0 U3201 ( .INP(n380), .ZN(n3810) );
  NAND2X1 U3202 ( .IN1(n2963), .IN2(n966), .QN(n2860) );
  INVX0 U3203 ( .INP(n314), .ZN(n3844) );
  INVX0 U3204 ( .INP(n315), .ZN(n3843) );
  INVX0 U3205 ( .INP(n316), .ZN(n3842) );
  INVX0 U3206 ( .INP(n317), .ZN(n3841) );
  INVX0 U3207 ( .INP(n318), .ZN(n3840) );
  INVX0 U3208 ( .INP(n319), .ZN(n3839) );
  INVX0 U3209 ( .INP(n320), .ZN(n3838) );
  INVX0 U3210 ( .INP(n321), .ZN(n3837) );
  INVX0 U3211 ( .INP(n322), .ZN(n3836) );
  INVX0 U3212 ( .INP(n323), .ZN(n3835) );
  INVX0 U3213 ( .INP(n324), .ZN(n3834) );
  INVX0 U3214 ( .INP(n325), .ZN(n3833) );
  INVX0 U3215 ( .INP(n326), .ZN(n3832) );
  INVX0 U3216 ( .INP(n327), .ZN(n3831) );
  INVX0 U3217 ( .INP(n328), .ZN(n3830) );
  INVX0 U3218 ( .INP(n329), .ZN(n3829) );
  INVX0 U3219 ( .INP(n330), .ZN(n3828) );
  INVX0 U3220 ( .INP(n331), .ZN(n3827) );
  INVX0 U3221 ( .INP(n332), .ZN(n3826) );
  INVX0 U3222 ( .INP(n333), .ZN(n3825) );
  INVX0 U3223 ( .INP(n334), .ZN(n3824) );
  INVX0 U3224 ( .INP(n335), .ZN(n3823) );
  INVX0 U3225 ( .INP(n336), .ZN(n3822) );
  INVX0 U3226 ( .INP(n337), .ZN(n3821) );
  INVX0 U3227 ( .INP(n338), .ZN(n3820) );
  INVX0 U3228 ( .INP(n339), .ZN(n3819) );
  INVX0 U3229 ( .INP(n340), .ZN(n3818) );
  INVX0 U3230 ( .INP(n341), .ZN(n3817) );
  INVX0 U3231 ( .INP(n342), .ZN(n3816) );
  INVX0 U3232 ( .INP(n343), .ZN(n3815) );
  NOR2X0 U3233 ( .IN1(n3489), .IN2(n3840), .QN(n2946) );
  INVX0 U3234 ( .INP(n313), .ZN(n3845) );
  NOR2X0 U3235 ( .IN1(n972), .IN2(n3223), .QN(n2965) );
  NOR2X0 U3236 ( .IN1(n3489), .IN2(n3844), .QN(n2958) );
  NOR2X0 U3237 ( .IN1(n3489), .IN2(n3843), .QN(n2955) );
  NOR2X0 U3238 ( .IN1(n3489), .IN2(n3842), .QN(n2952) );
  NOR2X0 U3239 ( .IN1(n3489), .IN2(n3841), .QN(n2949) );
  NOR2X0 U3240 ( .IN1(n3849), .IN2(N18), .QN(n2812) );
  NOR2X0 U3241 ( .IN1(n3853), .IN2(N22), .QN(n2500) );
  NOR2X0 U3242 ( .IN1(n3848), .IN2(N17), .QN(n2815) );
  NOR2X0 U3243 ( .IN1(n3852), .IN2(N21), .QN(n2503) );
  NOR2X0 U3244 ( .IN1(n3847), .IN2(N20), .QN(n2818) );
  NOR2X0 U3245 ( .IN1(n3851), .IN2(N24), .QN(n2506) );
  NOR2X0 U3246 ( .IN1(n3846), .IN2(N19), .QN(n2820) );
  NOR2X0 U3247 ( .IN1(n3850), .IN2(N23), .QN(n2508) );
  NOR2X0 U3248 ( .IN1(N17), .IN2(N18), .QN(n2814) );
  NOR2X0 U3249 ( .IN1(N21), .IN2(N22), .QN(n2502) );
  NOR2X0 U3250 ( .IN1(N19), .IN2(N20), .QN(n2813) );
  NOR2X0 U3251 ( .IN1(N23), .IN2(N24), .QN(n2501) );
  INVX0 U3252 ( .INP(N17), .ZN(n3849) );
  INVX0 U3253 ( .INP(N21), .ZN(n3853) );
  INVX0 U3254 ( .INP(N19), .ZN(n3847) );
  INVX0 U3255 ( .INP(N23), .ZN(n3851) );
  INVX0 U3256 ( .INP(N18), .ZN(n3848) );
  INVX0 U3257 ( .INP(N20), .ZN(n3846) );
  INVX0 U3258 ( .INP(N22), .ZN(n3852) );
  INVX0 U3259 ( .INP(N24), .ZN(n3850) );
  INVX0 U3260 ( .INP(rst), .ZN(n3772) );
  INVX0 U3261 ( .INP(rst), .ZN(n3776) );
  INVX0 U3262 ( .INP(rst), .ZN(n3775) );
  INVX0 U3263 ( .INP(rst), .ZN(n3774) );
  INVX0 U3264 ( .INP(rst), .ZN(n3773) );
  INVX0 U3265 ( .INP(rst), .ZN(n3771) );
  INVX0 U3266 ( .INP(rst), .ZN(n3770) );
  INVX0 U3267 ( .INP(rst), .ZN(n3777) );
  NBUFFX2 U3268 ( .INP(n3812), .Z(n3484) );
  NBUFFX2 U3269 ( .INP(n3812), .Z(n3485) );
  NBUFFX2 U3270 ( .INP(n3813), .Z(n3487) );
  NBUFFX2 U3271 ( .INP(n2867), .Z(n3492) );
  NBUFFX2 U3272 ( .INP(n2867), .Z(n3493) );
  NBUFFX2 U3273 ( .INP(n2867), .Z(n3494) );
  NBUFFX2 U3274 ( .INP(n2863), .Z(n3495) );
  NBUFFX2 U3275 ( .INP(n2863), .Z(n3496) );
  NBUFFX2 U3276 ( .INP(n2863), .Z(n3497) );
  NBUFFX2 U3277 ( .INP(n2863), .Z(n3498) );
  NBUFFX2 U3278 ( .INP(n2863), .Z(n3499) );
  NBUFFX2 U3279 ( .INP(n2535), .Z(n3628) );
  NBUFFX2 U3280 ( .INP(n2535), .Z(n3629) );
  NBUFFX2 U3281 ( .INP(n2534), .Z(n3631) );
  NBUFFX2 U3282 ( .INP(n2534), .Z(n3632) );
  NBUFFX2 U3283 ( .INP(n2532), .Z(n3634) );
  NBUFFX2 U3284 ( .INP(n2532), .Z(n3635) );
  NBUFFX2 U3285 ( .INP(n2531), .Z(n3637) );
  NBUFFX2 U3286 ( .INP(n2531), .Z(n3638) );
  NBUFFX2 U3287 ( .INP(n2530), .Z(n3640) );
  NBUFFX2 U3288 ( .INP(n2530), .Z(n3641) );
  NBUFFX2 U3289 ( .INP(n2529), .Z(n3643) );
  NBUFFX2 U3290 ( .INP(n2529), .Z(n3644) );
  NBUFFX2 U3291 ( .INP(n2527), .Z(n3646) );
  NBUFFX2 U3292 ( .INP(n2527), .Z(n3647) );
  NBUFFX2 U3293 ( .INP(n2526), .Z(n3649) );
  NBUFFX2 U3294 ( .INP(n2526), .Z(n3650) );
  NBUFFX2 U3295 ( .INP(n2525), .Z(n3652) );
  NBUFFX2 U3296 ( .INP(n2525), .Z(n3653) );
  NBUFFX2 U3297 ( .INP(n2524), .Z(n3655) );
  NBUFFX2 U3298 ( .INP(n2524), .Z(n3656) );
  NBUFFX2 U3299 ( .INP(n2522), .Z(n3658) );
  NBUFFX2 U3300 ( .INP(n2522), .Z(n3659) );
  NBUFFX2 U3301 ( .INP(n2521), .Z(n3661) );
  NBUFFX2 U3302 ( .INP(n2521), .Z(n3662) );
  NBUFFX2 U3303 ( .INP(n2520), .Z(n3664) );
  NBUFFX2 U3304 ( .INP(n2520), .Z(n3665) );
  NBUFFX2 U3305 ( .INP(n2519), .Z(n3667) );
  NBUFFX2 U3306 ( .INP(n2519), .Z(n3668) );
  NBUFFX2 U3307 ( .INP(n2517), .Z(n3670) );
  NBUFFX2 U3308 ( .INP(n2517), .Z(n3671) );
  NBUFFX2 U3309 ( .INP(n2516), .Z(n3673) );
  NBUFFX2 U3310 ( .INP(n2516), .Z(n3674) );
  NBUFFX2 U3311 ( .INP(n2223), .Z(n3676) );
  NBUFFX2 U3312 ( .INP(n2223), .Z(n3677) );
  NBUFFX2 U3313 ( .INP(n2222), .Z(n3679) );
  NBUFFX2 U3314 ( .INP(n2222), .Z(n3680) );
  NBUFFX2 U3315 ( .INP(n2220), .Z(n3682) );
  NBUFFX2 U3316 ( .INP(n2220), .Z(n3683) );
  NBUFFX2 U3317 ( .INP(n2219), .Z(n3685) );
  NBUFFX2 U3318 ( .INP(n2219), .Z(n3686) );
  NBUFFX2 U3319 ( .INP(n2218), .Z(n3688) );
  NBUFFX2 U3320 ( .INP(n2218), .Z(n3689) );
  NBUFFX2 U3321 ( .INP(n2217), .Z(n3691) );
  NBUFFX2 U3322 ( .INP(n2217), .Z(n3692) );
  NBUFFX2 U3323 ( .INP(n2215), .Z(n3694) );
  NBUFFX2 U3324 ( .INP(n2215), .Z(n3695) );
  NBUFFX2 U3325 ( .INP(n2214), .Z(n3697) );
  NBUFFX2 U3326 ( .INP(n2214), .Z(n3698) );
  NBUFFX2 U3327 ( .INP(n2213), .Z(n3700) );
  NBUFFX2 U3328 ( .INP(n2213), .Z(n3701) );
  NBUFFX2 U3329 ( .INP(n2212), .Z(n3703) );
  NBUFFX2 U3330 ( .INP(n2212), .Z(n3704) );
  NBUFFX2 U3331 ( .INP(n2210), .Z(n3706) );
  NBUFFX2 U3332 ( .INP(n2210), .Z(n3707) );
  NBUFFX2 U3333 ( .INP(n2209), .Z(n3709) );
  NBUFFX2 U3334 ( .INP(n2209), .Z(n3710) );
  NBUFFX2 U3335 ( .INP(n2208), .Z(n3712) );
  NBUFFX2 U3336 ( .INP(n2208), .Z(n3713) );
  NBUFFX2 U3337 ( .INP(n2207), .Z(n3715) );
  NBUFFX2 U3338 ( .INP(n2207), .Z(n3716) );
  NBUFFX2 U3339 ( .INP(n2205), .Z(n3718) );
  NBUFFX2 U3340 ( .INP(n2205), .Z(n3719) );
  NBUFFX2 U3341 ( .INP(n2204), .Z(n3721) );
  NBUFFX2 U3342 ( .INP(n2204), .Z(n3722) );
  INVX0 U3343 ( .INP(n3483), .ZN(n3491) );
  INVX0 U3344 ( .INP(n3500), .ZN(n3507) );
  INVX0 U3345 ( .INP(n3508), .ZN(n3515) );
  INVX0 U3346 ( .INP(n3516), .ZN(n3523) );
  INVX0 U3347 ( .INP(n3524), .ZN(n3531) );
  INVX0 U3348 ( .INP(n3532), .ZN(n3539) );
  INVX0 U3349 ( .INP(n3540), .ZN(n3547) );
  INVX0 U3350 ( .INP(n3548), .ZN(n3555) );
  INVX0 U3351 ( .INP(n3556), .ZN(n3563) );
  INVX0 U3352 ( .INP(n3564), .ZN(n3571) );
  INVX0 U3353 ( .INP(n3572), .ZN(n3579) );
  INVX0 U3354 ( .INP(n3580), .ZN(n3587) );
  INVX0 U3355 ( .INP(n3588), .ZN(n3595) );
  INVX0 U3356 ( .INP(n3596), .ZN(n3603) );
  INVX0 U3357 ( .INP(n3604), .ZN(n3611) );
  INVX0 U3358 ( .INP(n3612), .ZN(n3619) );
  INVX0 U3359 ( .INP(n3620), .ZN(n3627) );
  INVX0 U3360 ( .INP(n3772), .ZN(n3724) );
  INVX0 U3361 ( .INP(n3772), .ZN(n3725) );
  INVX0 U3362 ( .INP(n3772), .ZN(n3726) );
  INVX0 U3363 ( .INP(n3772), .ZN(n3727) );
  INVX0 U3364 ( .INP(n3772), .ZN(n3728) );
  INVX0 U3365 ( .INP(n3772), .ZN(n3729) );
  INVX0 U3366 ( .INP(n3772), .ZN(n3730) );
  INVX0 U3367 ( .INP(n3772), .ZN(n3731) );
  INVX0 U3368 ( .INP(n3772), .ZN(n3732) );
  INVX0 U3369 ( .INP(n3771), .ZN(n3733) );
  INVX0 U3370 ( .INP(n3771), .ZN(n3734) );
  INVX0 U3371 ( .INP(n3771), .ZN(n3735) );
  INVX0 U3372 ( .INP(n3771), .ZN(n3736) );
  INVX0 U3373 ( .INP(n3771), .ZN(n3737) );
  INVX0 U3374 ( .INP(n3771), .ZN(n3738) );
  INVX0 U3375 ( .INP(n3771), .ZN(n3739) );
  INVX0 U3376 ( .INP(n3771), .ZN(n3740) );
  INVX0 U3377 ( .INP(n3771), .ZN(n3741) );
  INVX0 U3378 ( .INP(n3771), .ZN(n3742) );
  INVX0 U3379 ( .INP(n3771), .ZN(n3743) );
  INVX0 U3380 ( .INP(n3771), .ZN(n3744) );
  INVX0 U3381 ( .INP(n3770), .ZN(n3745) );
  INVX0 U3382 ( .INP(n3770), .ZN(n3746) );
  INVX0 U3383 ( .INP(n3770), .ZN(n3747) );
  INVX0 U3384 ( .INP(n3770), .ZN(n3748) );
  INVX0 U3385 ( .INP(n3770), .ZN(n3749) );
  INVX0 U3386 ( .INP(n3770), .ZN(n3750) );
  INVX0 U3387 ( .INP(n3770), .ZN(n3751) );
  INVX0 U3388 ( .INP(n3770), .ZN(n3752) );
  INVX0 U3389 ( .INP(n3770), .ZN(n3753) );
  INVX0 U3390 ( .INP(n3770), .ZN(n3754) );
  INVX0 U3391 ( .INP(n3770), .ZN(n3755) );
  INVX0 U3392 ( .INP(n3770), .ZN(n3756) );
  INVX0 U3393 ( .INP(n3769), .ZN(n3757) );
  INVX0 U3394 ( .INP(n3769), .ZN(n3758) );
  INVX0 U3395 ( .INP(n3769), .ZN(n3759) );
  INVX0 U3396 ( .INP(n3769), .ZN(n3760) );
  INVX0 U3397 ( .INP(n3769), .ZN(n3761) );
  INVX0 U3398 ( .INP(n3769), .ZN(n3762) );
  INVX0 U3399 ( .INP(n3769), .ZN(n3763) );
  INVX0 U3400 ( .INP(n3769), .ZN(n3764) );
endmodule



module thumb_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   \carry[1] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34;

  AND2X1 U1 ( .IN1(A[30]), .IN2(n2), .Q(n1) );
  AND2X1 U2 ( .IN1(A[29]), .IN2(n3), .Q(n2) );
  AND2X1 U3 ( .IN1(A[28]), .IN2(n4), .Q(n3) );
  AND2X1 U4 ( .IN1(A[27]), .IN2(n5), .Q(n4) );
  AND2X1 U5 ( .IN1(A[26]), .IN2(n6), .Q(n5) );
  AND2X1 U6 ( .IN1(A[25]), .IN2(n7), .Q(n6) );
  AND2X1 U7 ( .IN1(A[24]), .IN2(n8), .Q(n7) );
  AND2X1 U8 ( .IN1(A[23]), .IN2(n9), .Q(n8) );
  AND2X1 U9 ( .IN1(A[22]), .IN2(n10), .Q(n9) );
  AND2X1 U10 ( .IN1(A[21]), .IN2(n11), .Q(n10) );
  AND2X1 U11 ( .IN1(A[20]), .IN2(n12), .Q(n11) );
  AND2X1 U12 ( .IN1(A[19]), .IN2(n13), .Q(n12) );
  AND2X1 U13 ( .IN1(A[18]), .IN2(n14), .Q(n13) );
  AND2X1 U14 ( .IN1(A[17]), .IN2(n15), .Q(n14) );
  AND2X1 U15 ( .IN1(A[16]), .IN2(n16), .Q(n15) );
  AND2X1 U16 ( .IN1(A[15]), .IN2(n17), .Q(n16) );
  AND2X1 U17 ( .IN1(A[14]), .IN2(n18), .Q(n17) );
  AND2X1 U18 ( .IN1(A[13]), .IN2(n19), .Q(n18) );
  AND2X1 U19 ( .IN1(A[12]), .IN2(n20), .Q(n19) );
  AND2X1 U20 ( .IN1(A[11]), .IN2(n21), .Q(n20) );
  AND2X1 U21 ( .IN1(A[10]), .IN2(n22), .Q(n21) );
  AND2X1 U22 ( .IN1(A[9]), .IN2(n23), .Q(n22) );
  AND2X1 U23 ( .IN1(A[8]), .IN2(n24), .Q(n23) );
  AND2X1 U24 ( .IN1(A[7]), .IN2(n25), .Q(n24) );
  AND2X1 U25 ( .IN1(A[6]), .IN2(n26), .Q(n25) );
  AND2X1 U26 ( .IN1(A[5]), .IN2(n27), .Q(n26) );
  AND2X1 U27 ( .IN1(A[4]), .IN2(n28), .Q(n27) );
  AND2X1 U28 ( .IN1(A[3]), .IN2(n29), .Q(n28) );
  AND2X1 U29 ( .IN1(A[2]), .IN2(n31), .Q(n29) );
  AND2X1 U30 ( .IN1(A[31]), .IN2(n1), .Q(n30) );
  AND2X1 U31 ( .IN1(A[1]), .IN2(\carry[1] ), .Q(n31) );
  NAND2X1 U32 ( .IN1(n32), .IN2(n33), .QN(\carry[1] ) );
  INVX0 U33 ( .INP(A[0]), .ZN(n32) );
  INVX0 U34 ( .INP(n34), .ZN(n33) );
  INVX0 U35 ( .INP(B[0]), .ZN(n34) );
  XOR2X1 U36 ( .IN1(n33), .IN2(A[0]), .Q(SUM[0]) );
  XOR2X1 U37 ( .IN1(A[10]), .IN2(n22), .Q(SUM[10]) );
  XOR2X1 U38 ( .IN1(A[11]), .IN2(n21), .Q(SUM[11]) );
  XOR2X1 U39 ( .IN1(A[12]), .IN2(n20), .Q(SUM[12]) );
  XOR2X1 U40 ( .IN1(A[13]), .IN2(n19), .Q(SUM[13]) );
  XOR2X1 U41 ( .IN1(A[14]), .IN2(n18), .Q(SUM[14]) );
  XOR2X1 U42 ( .IN1(A[15]), .IN2(n17), .Q(SUM[15]) );
  XOR2X1 U43 ( .IN1(A[16]), .IN2(n16), .Q(SUM[16]) );
  XOR2X1 U44 ( .IN1(A[17]), .IN2(n15), .Q(SUM[17]) );
  XOR2X1 U45 ( .IN1(A[18]), .IN2(n14), .Q(SUM[18]) );
  XOR2X1 U46 ( .IN1(A[19]), .IN2(n13), .Q(SUM[19]) );
  XOR2X1 U47 ( .IN1(A[1]), .IN2(\carry[1] ), .Q(SUM[1]) );
  XOR2X1 U48 ( .IN1(A[20]), .IN2(n12), .Q(SUM[20]) );
  XOR2X1 U49 ( .IN1(A[21]), .IN2(n11), .Q(SUM[21]) );
  XOR2X1 U50 ( .IN1(A[22]), .IN2(n10), .Q(SUM[22]) );
  XOR2X1 U51 ( .IN1(A[23]), .IN2(n9), .Q(SUM[23]) );
  XOR2X1 U52 ( .IN1(A[24]), .IN2(n8), .Q(SUM[24]) );
  XOR2X1 U53 ( .IN1(A[25]), .IN2(n7), .Q(SUM[25]) );
  XOR2X1 U54 ( .IN1(A[26]), .IN2(n6), .Q(SUM[26]) );
  XOR2X1 U55 ( .IN1(A[27]), .IN2(n5), .Q(SUM[27]) );
  XOR2X1 U56 ( .IN1(A[28]), .IN2(n4), .Q(SUM[28]) );
  XOR2X1 U57 ( .IN1(A[29]), .IN2(n3), .Q(SUM[29]) );
  XOR2X1 U58 ( .IN1(A[2]), .IN2(n31), .Q(SUM[2]) );
  XOR2X1 U59 ( .IN1(A[30]), .IN2(n2), .Q(SUM[30]) );
  XOR2X1 U60 ( .IN1(A[31]), .IN2(n1), .Q(SUM[31]) );
  XOR2X1 U61 ( .IN1(A[32]), .IN2(n30), .Q(SUM[32]) );
  XOR2X1 U62 ( .IN1(A[3]), .IN2(n29), .Q(SUM[3]) );
  XOR2X1 U63 ( .IN1(A[4]), .IN2(n28), .Q(SUM[4]) );
  XOR2X1 U64 ( .IN1(A[5]), .IN2(n27), .Q(SUM[5]) );
  XOR2X1 U65 ( .IN1(A[6]), .IN2(n26), .Q(SUM[6]) );
  XOR2X1 U66 ( .IN1(A[7]), .IN2(n25), .Q(SUM[7]) );
  XOR2X1 U67 ( .IN1(A[8]), .IN2(n24), .Q(SUM[8]) );
  XOR2X1 U68 ( .IN1(A[9]), .IN2(n23), .Q(SUM[9]) );
endmodule


module thumb_DW01_addsub_1 ( A, B, CI, ADD_SUB, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [33:0] carry;
  wire   [32:0] B_AS;

  FADDX1 U1_31 ( .A(A[31]), .B(B_AS[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B_AS[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B_AS[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B_AS[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B_AS[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B_AS[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B_AS[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B_AS[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B_AS[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B_AS[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B_AS[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B_AS[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B_AS[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B_AS[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B_AS[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B_AS[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B_AS[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FADDX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FADDX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FADDX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FADDX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FADDX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FADDX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FADDX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FADDX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0]) );
  XOR2X1 U1 ( .IN1(B_AS[32]), .IN2(carry[32]), .Q(SUM[32]) );
  XOR2X1 U2 ( .IN1(CI), .IN2(ADD_SUB), .Q(carry[0]) );
  XOR2X1 U3 ( .IN1(B[9]), .IN2(ADD_SUB), .Q(B_AS[9]) );
  XOR2X1 U4 ( .IN1(B[8]), .IN2(ADD_SUB), .Q(B_AS[8]) );
  XOR2X1 U5 ( .IN1(B[7]), .IN2(ADD_SUB), .Q(B_AS[7]) );
  XOR2X1 U6 ( .IN1(B[6]), .IN2(ADD_SUB), .Q(B_AS[6]) );
  XOR2X1 U7 ( .IN1(B[5]), .IN2(ADD_SUB), .Q(B_AS[5]) );
  XOR2X1 U8 ( .IN1(B[4]), .IN2(ADD_SUB), .Q(B_AS[4]) );
  XOR2X1 U9 ( .IN1(B[3]), .IN2(ADD_SUB), .Q(B_AS[3]) );
  XOR2X1 U10 ( .IN1(B[32]), .IN2(ADD_SUB), .Q(B_AS[32]) );
  XOR2X1 U11 ( .IN1(B[31]), .IN2(ADD_SUB), .Q(B_AS[31]) );
  XOR2X1 U12 ( .IN1(B[30]), .IN2(ADD_SUB), .Q(B_AS[30]) );
  XOR2X1 U13 ( .IN1(B[2]), .IN2(ADD_SUB), .Q(B_AS[2]) );
  XOR2X1 U14 ( .IN1(B[29]), .IN2(ADD_SUB), .Q(B_AS[29]) );
  XOR2X1 U15 ( .IN1(B[28]), .IN2(ADD_SUB), .Q(B_AS[28]) );
  XOR2X1 U16 ( .IN1(B[27]), .IN2(ADD_SUB), .Q(B_AS[27]) );
  XOR2X1 U17 ( .IN1(B[26]), .IN2(ADD_SUB), .Q(B_AS[26]) );
  XOR2X1 U18 ( .IN1(B[25]), .IN2(ADD_SUB), .Q(B_AS[25]) );
  XOR2X1 U19 ( .IN1(B[24]), .IN2(ADD_SUB), .Q(B_AS[24]) );
  XOR2X1 U20 ( .IN1(B[23]), .IN2(ADD_SUB), .Q(B_AS[23]) );
  XOR2X1 U21 ( .IN1(B[22]), .IN2(ADD_SUB), .Q(B_AS[22]) );
  XOR2X1 U22 ( .IN1(B[21]), .IN2(ADD_SUB), .Q(B_AS[21]) );
  XOR2X1 U23 ( .IN1(B[20]), .IN2(ADD_SUB), .Q(B_AS[20]) );
  XOR2X1 U24 ( .IN1(B[1]), .IN2(ADD_SUB), .Q(B_AS[1]) );
  XOR2X1 U25 ( .IN1(B[19]), .IN2(ADD_SUB), .Q(B_AS[19]) );
  XOR2X1 U26 ( .IN1(B[18]), .IN2(ADD_SUB), .Q(B_AS[18]) );
  XOR2X1 U27 ( .IN1(B[17]), .IN2(ADD_SUB), .Q(B_AS[17]) );
  XOR2X1 U28 ( .IN1(B[16]), .IN2(ADD_SUB), .Q(B_AS[16]) );
  XOR2X1 U29 ( .IN1(B[15]), .IN2(ADD_SUB), .Q(B_AS[15]) );
  XOR2X1 U30 ( .IN1(B[14]), .IN2(ADD_SUB), .Q(B_AS[14]) );
  XOR2X1 U31 ( .IN1(B[13]), .IN2(ADD_SUB), .Q(B_AS[13]) );
  XOR2X1 U32 ( .IN1(B[12]), .IN2(ADD_SUB), .Q(B_AS[12]) );
  XOR2X1 U33 ( .IN1(B[11]), .IN2(ADD_SUB), .Q(B_AS[11]) );
  XOR2X1 U34 ( .IN1(B[10]), .IN2(ADD_SUB), .Q(B_AS[10]) );
  XOR2X1 U35 ( .IN1(B[0]), .IN2(ADD_SUB), .Q(B_AS[0]) );
endmodule


module thumb_DW01_addsub_2 ( A, B, CI, ADD_SUB, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [33:0] carry;
  wire   [32:0] B_AS;
  assign carry[0] = ADD_SUB;

  FADDX1 U1_31 ( .A(A[31]), .B(carry[0]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(carry[0]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(carry[0]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(carry[0]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(carry[0]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(carry[0]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(carry[0]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(carry[0]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(carry[0]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(carry[0]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(carry[0]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(carry[0]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(carry[0]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(carry[0]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(carry[0]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(carry[0]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(carry[0]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(carry[0]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(carry[0]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(carry[0]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FADDX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FADDX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FADDX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FADDX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FADDX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FADDX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FADDX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FADDX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0]) );
  XOR2X1 U1 ( .IN1(carry[0]), .IN2(carry[32]), .Q(SUM[32]) );
  XOR2X1 U2 ( .IN1(B[9]), .IN2(carry[0]), .Q(B_AS[9]) );
  XOR2X1 U3 ( .IN1(B[8]), .IN2(carry[0]), .Q(B_AS[8]) );
  XOR2X1 U4 ( .IN1(B[7]), .IN2(carry[0]), .Q(B_AS[7]) );
  XOR2X1 U5 ( .IN1(B[6]), .IN2(carry[0]), .Q(B_AS[6]) );
  XOR2X1 U6 ( .IN1(B[5]), .IN2(carry[0]), .Q(B_AS[5]) );
  XOR2X1 U7 ( .IN1(B[4]), .IN2(carry[0]), .Q(B_AS[4]) );
  XOR2X1 U8 ( .IN1(B[3]), .IN2(carry[0]), .Q(B_AS[3]) );
  XOR2X1 U9 ( .IN1(B[2]), .IN2(carry[0]), .Q(B_AS[2]) );
  XOR2X1 U10 ( .IN1(B[1]), .IN2(carry[0]), .Q(B_AS[1]) );
  XOR2X1 U11 ( .IN1(B[11]), .IN2(carry[0]), .Q(B_AS[11]) );
  XOR2X1 U12 ( .IN1(B[10]), .IN2(carry[0]), .Q(B_AS[10]) );
  XOR2X1 U13 ( .IN1(B[0]), .IN2(carry[0]), .Q(B_AS[0]) );
endmodule


module thumb_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [32:1] carry;
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  AND2X1 U1 ( .IN1(A[1]), .IN2(B[1]), .Q(n1) );
  AND2X1 U2 ( .IN1(A[6]), .IN2(carry[6]), .Q(n2) );
  AND2X1 U3 ( .IN1(A[7]), .IN2(n2), .Q(n3) );
  AND2X1 U4 ( .IN1(A[8]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(A[9]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(A[10]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(A[11]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(A[12]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(A[13]), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(A[14]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(A[15]), .IN2(n10), .Q(n11) );
  AND2X1 U12 ( .IN1(A[16]), .IN2(n11), .Q(n12) );
  AND2X1 U13 ( .IN1(A[17]), .IN2(n12), .Q(n13) );
  AND2X1 U14 ( .IN1(A[18]), .IN2(n13), .Q(n14) );
  AND2X1 U15 ( .IN1(A[19]), .IN2(n14), .Q(n15) );
  AND2X1 U16 ( .IN1(A[20]), .IN2(n15), .Q(n16) );
  AND2X1 U17 ( .IN1(A[21]), .IN2(n16), .Q(n17) );
  AND2X1 U18 ( .IN1(A[22]), .IN2(n17), .Q(n18) );
  AND2X1 U19 ( .IN1(A[23]), .IN2(n18), .Q(n19) );
  AND2X1 U20 ( .IN1(A[24]), .IN2(n19), .Q(n20) );
  AND2X1 U21 ( .IN1(A[25]), .IN2(n20), .Q(n21) );
  AND2X1 U22 ( .IN1(A[26]), .IN2(n21), .Q(n22) );
  AND2X1 U23 ( .IN1(A[27]), .IN2(n22), .Q(n23) );
  AND2X1 U24 ( .IN1(A[28]), .IN2(n23), .Q(n24) );
  AND2X1 U25 ( .IN1(A[29]), .IN2(n24), .Q(n25) );
  AND2X1 U26 ( .IN1(A[30]), .IN2(n25), .Q(n26) );
  AND2X1 U27 ( .IN1(A[31]), .IN2(n26), .Q(SUM[32]) );
  XOR2X1 U28 ( .IN1(A[31]), .IN2(n26), .Q(SUM[31]) );
  XOR2X1 U29 ( .IN1(A[30]), .IN2(n25), .Q(SUM[30]) );
  XOR2X1 U30 ( .IN1(A[29]), .IN2(n24), .Q(SUM[29]) );
  XOR2X1 U31 ( .IN1(A[28]), .IN2(n23), .Q(SUM[28]) );
  XOR2X1 U32 ( .IN1(A[27]), .IN2(n22), .Q(SUM[27]) );
  XOR2X1 U33 ( .IN1(A[26]), .IN2(n21), .Q(SUM[26]) );
  XOR2X1 U34 ( .IN1(A[25]), .IN2(n20), .Q(SUM[25]) );
  XOR2X1 U35 ( .IN1(A[24]), .IN2(n19), .Q(SUM[24]) );
  XOR2X1 U36 ( .IN1(A[23]), .IN2(n18), .Q(SUM[23]) );
  XOR2X1 U37 ( .IN1(A[22]), .IN2(n17), .Q(SUM[22]) );
  XOR2X1 U38 ( .IN1(A[21]), .IN2(n16), .Q(SUM[21]) );
  XOR2X1 U39 ( .IN1(A[20]), .IN2(n15), .Q(SUM[20]) );
  XOR2X1 U40 ( .IN1(A[19]), .IN2(n14), .Q(SUM[19]) );
  XOR2X1 U41 ( .IN1(A[18]), .IN2(n13), .Q(SUM[18]) );
  XOR2X1 U42 ( .IN1(A[17]), .IN2(n12), .Q(SUM[17]) );
  XOR2X1 U43 ( .IN1(A[16]), .IN2(n11), .Q(SUM[16]) );
  XOR2X1 U44 ( .IN1(A[15]), .IN2(n10), .Q(SUM[15]) );
  XOR2X1 U45 ( .IN1(A[14]), .IN2(n9), .Q(SUM[14]) );
  XOR2X1 U46 ( .IN1(A[13]), .IN2(n8), .Q(SUM[13]) );
  XOR2X1 U47 ( .IN1(A[12]), .IN2(n7), .Q(SUM[12]) );
  XOR2X1 U48 ( .IN1(A[11]), .IN2(n6), .Q(SUM[11]) );
  XOR2X1 U49 ( .IN1(A[10]), .IN2(n5), .Q(SUM[10]) );
  XOR2X1 U50 ( .IN1(A[9]), .IN2(n4), .Q(SUM[9]) );
  XOR2X1 U51 ( .IN1(A[8]), .IN2(n3), .Q(SUM[8]) );
  XOR2X1 U52 ( .IN1(A[7]), .IN2(n2), .Q(SUM[7]) );
  XOR2X1 U53 ( .IN1(A[6]), .IN2(carry[6]), .Q(SUM[6]) );
  XOR2X1 U54 ( .IN1(A[1]), .IN2(B[1]), .Q(SUM[1]) );
endmodule


module thumb_DW01_add_1 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [32:1] carry;

  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(A[31]), .IN2(n28), .Q(SUM[32]) );
  AND2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(n2) );
  AND2X1 U3 ( .IN1(A[5]), .IN2(carry[5]), .Q(n3) );
  AND2X1 U4 ( .IN1(A[6]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(A[7]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(A[8]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(A[9]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(A[10]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(A[11]), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(A[12]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(A[13]), .IN2(n10), .Q(n11) );
  AND2X1 U12 ( .IN1(A[14]), .IN2(n11), .Q(n12) );
  AND2X1 U13 ( .IN1(A[15]), .IN2(n12), .Q(n13) );
  AND2X1 U14 ( .IN1(A[16]), .IN2(n13), .Q(n14) );
  AND2X1 U15 ( .IN1(A[17]), .IN2(n14), .Q(n15) );
  AND2X1 U16 ( .IN1(A[18]), .IN2(n15), .Q(n16) );
  AND2X1 U17 ( .IN1(A[19]), .IN2(n16), .Q(n17) );
  AND2X1 U18 ( .IN1(A[20]), .IN2(n17), .Q(n18) );
  AND2X1 U19 ( .IN1(A[21]), .IN2(n18), .Q(n19) );
  AND2X1 U20 ( .IN1(A[22]), .IN2(n19), .Q(n20) );
  AND2X1 U21 ( .IN1(A[23]), .IN2(n20), .Q(n21) );
  AND2X1 U22 ( .IN1(A[24]), .IN2(n21), .Q(n22) );
  AND2X1 U23 ( .IN1(A[25]), .IN2(n22), .Q(n23) );
  AND2X1 U24 ( .IN1(A[26]), .IN2(n23), .Q(n24) );
  AND2X1 U25 ( .IN1(A[27]), .IN2(n24), .Q(n25) );
  AND2X1 U26 ( .IN1(A[28]), .IN2(n25), .Q(n26) );
  AND2X1 U27 ( .IN1(A[29]), .IN2(n26), .Q(n27) );
  AND2X1 U28 ( .IN1(A[30]), .IN2(n27), .Q(n28) );
  XOR2X1 U29 ( .IN1(A[31]), .IN2(n28), .Q(SUM[31]) );
  XOR2X1 U30 ( .IN1(A[30]), .IN2(n27), .Q(SUM[30]) );
  XOR2X1 U31 ( .IN1(A[29]), .IN2(n26), .Q(SUM[29]) );
  XOR2X1 U32 ( .IN1(A[28]), .IN2(n25), .Q(SUM[28]) );
  XOR2X1 U33 ( .IN1(A[27]), .IN2(n24), .Q(SUM[27]) );
  XOR2X1 U34 ( .IN1(A[26]), .IN2(n23), .Q(SUM[26]) );
  XOR2X1 U35 ( .IN1(A[25]), .IN2(n22), .Q(SUM[25]) );
  XOR2X1 U36 ( .IN1(A[24]), .IN2(n21), .Q(SUM[24]) );
  XOR2X1 U37 ( .IN1(A[23]), .IN2(n20), .Q(SUM[23]) );
  XOR2X1 U38 ( .IN1(A[22]), .IN2(n19), .Q(SUM[22]) );
  XOR2X1 U39 ( .IN1(A[21]), .IN2(n18), .Q(SUM[21]) );
  XOR2X1 U40 ( .IN1(A[20]), .IN2(n17), .Q(SUM[20]) );
  XOR2X1 U41 ( .IN1(A[19]), .IN2(n16), .Q(SUM[19]) );
  XOR2X1 U42 ( .IN1(A[18]), .IN2(n15), .Q(SUM[18]) );
  XOR2X1 U43 ( .IN1(A[17]), .IN2(n14), .Q(SUM[17]) );
  XOR2X1 U44 ( .IN1(A[16]), .IN2(n13), .Q(SUM[16]) );
  XOR2X1 U45 ( .IN1(A[15]), .IN2(n12), .Q(SUM[15]) );
  XOR2X1 U46 ( .IN1(A[14]), .IN2(n11), .Q(SUM[14]) );
  XOR2X1 U47 ( .IN1(A[13]), .IN2(n10), .Q(SUM[13]) );
  XOR2X1 U48 ( .IN1(A[12]), .IN2(n9), .Q(SUM[12]) );
  XOR2X1 U49 ( .IN1(A[11]), .IN2(n8), .Q(SUM[11]) );
  XOR2X1 U50 ( .IN1(A[10]), .IN2(n7), .Q(SUM[10]) );
  XOR2X1 U51 ( .IN1(A[9]), .IN2(n6), .Q(SUM[9]) );
  XOR2X1 U52 ( .IN1(A[8]), .IN2(n5), .Q(SUM[8]) );
  XOR2X1 U53 ( .IN1(A[7]), .IN2(n4), .Q(SUM[7]) );
  XOR2X1 U54 ( .IN1(A[6]), .IN2(n3), .Q(SUM[6]) );
  XOR2X1 U55 ( .IN1(A[5]), .IN2(carry[5]), .Q(SUM[5]) );
  XOR2X1 U56 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module thumb_DW01_add_2 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [32:1] carry;
  assign SUM[1] = A[1];
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  AND2X1 U1 ( .IN1(A[2]), .IN2(B[2]), .Q(n1) );
  AND2X1 U2 ( .IN1(A[7]), .IN2(carry[7]), .Q(n2) );
  AND2X1 U3 ( .IN1(A[8]), .IN2(n2), .Q(n3) );
  AND2X1 U4 ( .IN1(A[9]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(A[10]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(A[11]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(A[12]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(A[13]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(A[14]), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(A[15]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(A[16]), .IN2(n10), .Q(n11) );
  AND2X1 U12 ( .IN1(A[17]), .IN2(n11), .Q(n12) );
  AND2X1 U13 ( .IN1(A[18]), .IN2(n12), .Q(n13) );
  AND2X1 U14 ( .IN1(A[19]), .IN2(n13), .Q(n14) );
  AND2X1 U15 ( .IN1(A[20]), .IN2(n14), .Q(n15) );
  AND2X1 U16 ( .IN1(A[21]), .IN2(n15), .Q(n16) );
  AND2X1 U17 ( .IN1(A[22]), .IN2(n16), .Q(n17) );
  AND2X1 U18 ( .IN1(A[23]), .IN2(n17), .Q(n18) );
  AND2X1 U19 ( .IN1(A[24]), .IN2(n18), .Q(n19) );
  AND2X1 U20 ( .IN1(A[25]), .IN2(n19), .Q(n20) );
  AND2X1 U21 ( .IN1(A[26]), .IN2(n20), .Q(n21) );
  AND2X1 U22 ( .IN1(A[27]), .IN2(n21), .Q(n22) );
  AND2X1 U23 ( .IN1(A[28]), .IN2(n22), .Q(n23) );
  AND2X1 U24 ( .IN1(A[29]), .IN2(n23), .Q(n24) );
  AND2X1 U25 ( .IN1(A[30]), .IN2(n24), .Q(n25) );
  AND2X1 U26 ( .IN1(A[31]), .IN2(n25), .Q(SUM[32]) );
  XOR2X1 U27 ( .IN1(A[31]), .IN2(n25), .Q(SUM[31]) );
  XOR2X1 U28 ( .IN1(A[30]), .IN2(n24), .Q(SUM[30]) );
  XOR2X1 U29 ( .IN1(A[29]), .IN2(n23), .Q(SUM[29]) );
  XOR2X1 U30 ( .IN1(A[28]), .IN2(n22), .Q(SUM[28]) );
  XOR2X1 U31 ( .IN1(A[27]), .IN2(n21), .Q(SUM[27]) );
  XOR2X1 U32 ( .IN1(A[26]), .IN2(n20), .Q(SUM[26]) );
  XOR2X1 U33 ( .IN1(A[25]), .IN2(n19), .Q(SUM[25]) );
  XOR2X1 U34 ( .IN1(A[24]), .IN2(n18), .Q(SUM[24]) );
  XOR2X1 U35 ( .IN1(A[23]), .IN2(n17), .Q(SUM[23]) );
  XOR2X1 U36 ( .IN1(A[22]), .IN2(n16), .Q(SUM[22]) );
  XOR2X1 U37 ( .IN1(A[21]), .IN2(n15), .Q(SUM[21]) );
  XOR2X1 U38 ( .IN1(A[20]), .IN2(n14), .Q(SUM[20]) );
  XOR2X1 U39 ( .IN1(A[19]), .IN2(n13), .Q(SUM[19]) );
  XOR2X1 U40 ( .IN1(A[18]), .IN2(n12), .Q(SUM[18]) );
  XOR2X1 U41 ( .IN1(A[17]), .IN2(n11), .Q(SUM[17]) );
  XOR2X1 U42 ( .IN1(A[16]), .IN2(n10), .Q(SUM[16]) );
  XOR2X1 U43 ( .IN1(A[15]), .IN2(n9), .Q(SUM[15]) );
  XOR2X1 U44 ( .IN1(A[14]), .IN2(n8), .Q(SUM[14]) );
  XOR2X1 U45 ( .IN1(A[13]), .IN2(n7), .Q(SUM[13]) );
  XOR2X1 U46 ( .IN1(A[12]), .IN2(n6), .Q(SUM[12]) );
  XOR2X1 U47 ( .IN1(A[11]), .IN2(n5), .Q(SUM[11]) );
  XOR2X1 U48 ( .IN1(A[10]), .IN2(n4), .Q(SUM[10]) );
  XOR2X1 U49 ( .IN1(A[9]), .IN2(n3), .Q(SUM[9]) );
  XOR2X1 U50 ( .IN1(A[8]), .IN2(n2), .Q(SUM[8]) );
  XOR2X1 U51 ( .IN1(A[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U52 ( .IN1(A[2]), .IN2(B[2]), .Q(SUM[2]) );
endmodule


module thumb_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;
  wire   [33:0] carry;

  FADDX1 U2_31 ( .A(A[31]), .B(n35), .CI(carry[31]), .CO(carry[32]), .S(
        DIFF[31]) );
  FADDX1 U2_30 ( .A(A[30]), .B(n34), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  FADDX1 U2_29 ( .A(A[29]), .B(n33), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  FADDX1 U2_28 ( .A(A[28]), .B(n32), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  FADDX1 U2_27 ( .A(A[27]), .B(n31), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  FADDX1 U2_26 ( .A(A[26]), .B(n30), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  FADDX1 U2_25 ( .A(A[25]), .B(n29), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  FADDX1 U2_24 ( .A(A[24]), .B(n28), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  FADDX1 U2_23 ( .A(A[23]), .B(n27), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1 U2_22 ( .A(A[22]), .B(n26), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n25), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n24), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n23), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n22), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n21), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n20), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n19), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n18), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n17), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n16), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n15), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n14), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n13), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n12), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_7 ( .A(A[7]), .B(n11), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  FADDX1 U2_6 ( .A(A[6]), .B(n10), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FADDX1 U2_5 ( .A(A[5]), .B(n9), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n8), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n7), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1 U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FADDX1 U2_1 ( .A(A[1]), .B(n5), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INVX0 U1 ( .INP(carry[32]), .ZN(DIFF[32]) );
  INVX0 U2 ( .INP(n4), .ZN(n2) );
  INVX0 U3 ( .INP(B[0]), .ZN(n4) );
  INVX0 U4 ( .INP(B[3]), .ZN(n7) );
  INVX0 U5 ( .INP(B[4]), .ZN(n8) );
  INVX0 U6 ( .INP(B[2]), .ZN(n6) );
  INVX0 U7 ( .INP(B[5]), .ZN(n9) );
  INVX0 U8 ( .INP(B[6]), .ZN(n10) );
  INVX0 U9 ( .INP(B[7]), .ZN(n11) );
  INVX0 U10 ( .INP(B[8]), .ZN(n12) );
  INVX0 U11 ( .INP(B[9]), .ZN(n13) );
  INVX0 U12 ( .INP(B[10]), .ZN(n14) );
  INVX0 U13 ( .INP(B[11]), .ZN(n15) );
  INVX0 U14 ( .INP(B[12]), .ZN(n16) );
  INVX0 U15 ( .INP(B[13]), .ZN(n17) );
  INVX0 U16 ( .INP(B[14]), .ZN(n18) );
  INVX0 U17 ( .INP(B[15]), .ZN(n19) );
  INVX0 U18 ( .INP(B[16]), .ZN(n20) );
  INVX0 U19 ( .INP(B[17]), .ZN(n21) );
  INVX0 U20 ( .INP(B[18]), .ZN(n22) );
  INVX0 U21 ( .INP(B[19]), .ZN(n23) );
  INVX0 U22 ( .INP(B[20]), .ZN(n24) );
  INVX0 U23 ( .INP(B[21]), .ZN(n25) );
  INVX0 U24 ( .INP(B[22]), .ZN(n26) );
  INVX0 U25 ( .INP(B[23]), .ZN(n27) );
  INVX0 U26 ( .INP(B[24]), .ZN(n28) );
  INVX0 U27 ( .INP(B[25]), .ZN(n29) );
  INVX0 U28 ( .INP(B[26]), .ZN(n30) );
  INVX0 U29 ( .INP(B[27]), .ZN(n31) );
  INVX0 U30 ( .INP(B[28]), .ZN(n32) );
  INVX0 U31 ( .INP(B[29]), .ZN(n33) );
  INVX0 U32 ( .INP(B[30]), .ZN(n34) );
  NAND2X1 U33 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U34 ( .INP(B[1]), .ZN(n5) );
  INVX0 U35 ( .INP(A[0]), .ZN(n1) );
  INVX0 U36 ( .INP(B[31]), .ZN(n35) );
  XOR2X1 U37 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module thumb_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59;
  wire   [33:0] carry;

  FADDX1 U2_7 ( .A(A[7]), .B(n52), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  FADDX1 U2_6 ( .A(A[6]), .B(n53), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FADDX1 U2_5 ( .A(A[5]), .B(n54), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  FADDX1 U2_4 ( .A(A[4]), .B(n55), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  FADDX1 U2_3 ( .A(A[3]), .B(n56), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n57), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n58), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  INVX0 U1 ( .INP(A[30]), .ZN(n45) );
  INVX0 U2 ( .INP(A[29]), .ZN(n44) );
  INVX0 U3 ( .INP(A[28]), .ZN(n43) );
  INVX0 U4 ( .INP(A[27]), .ZN(n42) );
  INVX0 U5 ( .INP(A[26]), .ZN(n41) );
  INVX0 U6 ( .INP(A[25]), .ZN(n40) );
  INVX0 U7 ( .INP(A[24]), .ZN(n39) );
  INVX0 U8 ( .INP(A[23]), .ZN(n38) );
  INVX0 U9 ( .INP(A[22]), .ZN(n37) );
  INVX0 U10 ( .INP(A[21]), .ZN(n36) );
  INVX0 U11 ( .INP(A[20]), .ZN(n35) );
  INVX0 U12 ( .INP(A[19]), .ZN(n34) );
  INVX0 U13 ( .INP(A[18]), .ZN(n33) );
  INVX0 U14 ( .INP(A[17]), .ZN(n32) );
  INVX0 U15 ( .INP(A[16]), .ZN(n31) );
  INVX0 U16 ( .INP(A[15]), .ZN(n30) );
  INVX0 U17 ( .INP(A[14]), .ZN(n29) );
  INVX0 U18 ( .INP(A[13]), .ZN(n28) );
  INVX0 U19 ( .INP(A[12]), .ZN(n27) );
  INVX0 U20 ( .INP(A[11]), .ZN(n26) );
  INVX0 U21 ( .INP(A[10]), .ZN(n25) );
  INVX0 U22 ( .INP(A[9]), .ZN(n49) );
  INVX0 U23 ( .INP(A[8]), .ZN(n47) );
  INVX0 U24 ( .INP(A[31]), .ZN(n46) );
  INVX0 U25 ( .INP(carry[8]), .ZN(n48) );
  INVX0 U26 ( .INP(n59), .ZN(n51) );
  INVX0 U27 ( .INP(B[0]), .ZN(n59) );
  INVX0 U28 ( .INP(B[3]), .ZN(n56) );
  INVX0 U29 ( .INP(B[4]), .ZN(n55) );
  INVX0 U30 ( .INP(B[2]), .ZN(n57) );
  INVX0 U31 ( .INP(B[5]), .ZN(n54) );
  INVX0 U32 ( .INP(B[6]), .ZN(n53) );
  NAND2X1 U33 ( .IN1(n50), .IN2(n51), .QN(carry[1]) );
  INVX0 U34 ( .INP(B[1]), .ZN(n58) );
  INVX0 U35 ( .INP(A[0]), .ZN(n50) );
  INVX0 U36 ( .INP(B[7]), .ZN(n52) );
  AND2X1 U37 ( .IN1(n47), .IN2(n48), .Q(n1) );
  AND2X1 U38 ( .IN1(n49), .IN2(n1), .Q(n2) );
  AND2X1 U39 ( .IN1(n25), .IN2(n2), .Q(n3) );
  AND2X1 U40 ( .IN1(n26), .IN2(n3), .Q(n4) );
  AND2X1 U41 ( .IN1(n27), .IN2(n4), .Q(n5) );
  AND2X1 U42 ( .IN1(n28), .IN2(n5), .Q(n6) );
  AND2X1 U43 ( .IN1(n29), .IN2(n6), .Q(n7) );
  AND2X1 U44 ( .IN1(n30), .IN2(n7), .Q(n8) );
  AND2X1 U45 ( .IN1(n31), .IN2(n8), .Q(n9) );
  AND2X1 U46 ( .IN1(n32), .IN2(n9), .Q(n10) );
  AND2X1 U47 ( .IN1(n33), .IN2(n10), .Q(n11) );
  AND2X1 U48 ( .IN1(n34), .IN2(n11), .Q(n12) );
  AND2X1 U49 ( .IN1(n35), .IN2(n12), .Q(n13) );
  AND2X1 U50 ( .IN1(n36), .IN2(n13), .Q(n14) );
  AND2X1 U51 ( .IN1(n37), .IN2(n14), .Q(n15) );
  AND2X1 U52 ( .IN1(n38), .IN2(n15), .Q(n16) );
  AND2X1 U53 ( .IN1(n39), .IN2(n16), .Q(n17) );
  AND2X1 U54 ( .IN1(n40), .IN2(n17), .Q(n18) );
  AND2X1 U55 ( .IN1(n41), .IN2(n18), .Q(n19) );
  AND2X1 U56 ( .IN1(n42), .IN2(n19), .Q(n20) );
  AND2X1 U57 ( .IN1(n43), .IN2(n20), .Q(n21) );
  AND2X1 U58 ( .IN1(n44), .IN2(n21), .Q(n22) );
  AND2X1 U59 ( .IN1(n45), .IN2(n22), .Q(n23) );
  AND2X1 U60 ( .IN1(n46), .IN2(n23), .Q(DIFF[32]) );
  XOR2X1 U61 ( .IN1(n2), .IN2(A[10]), .Q(DIFF[10]) );
  XOR2X1 U62 ( .IN1(n3), .IN2(A[11]), .Q(DIFF[11]) );
  XOR2X1 U63 ( .IN1(n4), .IN2(A[12]), .Q(DIFF[12]) );
  XOR2X1 U64 ( .IN1(n5), .IN2(A[13]), .Q(DIFF[13]) );
  XOR2X1 U65 ( .IN1(n6), .IN2(A[14]), .Q(DIFF[14]) );
  XOR2X1 U66 ( .IN1(n7), .IN2(A[15]), .Q(DIFF[15]) );
  XOR2X1 U67 ( .IN1(n8), .IN2(A[16]), .Q(DIFF[16]) );
  XOR2X1 U68 ( .IN1(n9), .IN2(A[17]), .Q(DIFF[17]) );
  XOR2X1 U69 ( .IN1(n10), .IN2(A[18]), .Q(DIFF[18]) );
  XOR2X1 U70 ( .IN1(n11), .IN2(A[19]), .Q(DIFF[19]) );
  XOR2X1 U71 ( .IN1(n12), .IN2(A[20]), .Q(DIFF[20]) );
  XOR2X1 U72 ( .IN1(n13), .IN2(A[21]), .Q(DIFF[21]) );
  XOR2X1 U73 ( .IN1(n14), .IN2(A[22]), .Q(DIFF[22]) );
  XOR2X1 U74 ( .IN1(n15), .IN2(A[23]), .Q(DIFF[23]) );
  XOR2X1 U75 ( .IN1(n16), .IN2(A[24]), .Q(DIFF[24]) );
  XOR2X1 U76 ( .IN1(n17), .IN2(A[25]), .Q(DIFF[25]) );
  XOR2X1 U77 ( .IN1(n18), .IN2(A[26]), .Q(DIFF[26]) );
  XOR2X1 U78 ( .IN1(n19), .IN2(A[27]), .Q(DIFF[27]) );
  XOR2X1 U79 ( .IN1(n20), .IN2(A[28]), .Q(DIFF[28]) );
  XOR2X1 U80 ( .IN1(n21), .IN2(A[29]), .Q(DIFF[29]) );
  XOR2X1 U81 ( .IN1(n22), .IN2(A[30]), .Q(DIFF[30]) );
  XOR2X1 U82 ( .IN1(n23), .IN2(A[31]), .Q(DIFF[31]) );
  XOR2X1 U83 ( .IN1(n48), .IN2(A[8]), .Q(DIFF[8]) );
  XOR2X1 U84 ( .IN1(n1), .IN2(A[9]), .Q(DIFF[9]) );
  XOR2X1 U85 ( .IN1(n51), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module thumb_DW01_add_3 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22;
  wire   [32:1] carry;
  assign SUM[1] = A[1];
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  AND2X1 U1 ( .IN1(A[2]), .IN2(B[2]), .Q(n1) );
  AND2X1 U2 ( .IN1(A[10]), .IN2(carry[10]), .Q(n2) );
  AND2X1 U3 ( .IN1(A[11]), .IN2(n2), .Q(n3) );
  AND2X1 U4 ( .IN1(A[12]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(A[13]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(A[14]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(A[15]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(A[16]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(A[17]), .IN2(n8), .Q(n9) );
  AND2X1 U10 ( .IN1(A[18]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(A[19]), .IN2(n10), .Q(n11) );
  AND2X1 U12 ( .IN1(A[20]), .IN2(n11), .Q(n12) );
  AND2X1 U13 ( .IN1(A[21]), .IN2(n12), .Q(n13) );
  AND2X1 U14 ( .IN1(A[22]), .IN2(n13), .Q(n14) );
  AND2X1 U15 ( .IN1(A[23]), .IN2(n14), .Q(n15) );
  AND2X1 U16 ( .IN1(A[24]), .IN2(n15), .Q(n16) );
  AND2X1 U17 ( .IN1(A[25]), .IN2(n16), .Q(n17) );
  AND2X1 U18 ( .IN1(A[26]), .IN2(n17), .Q(n18) );
  AND2X1 U19 ( .IN1(A[27]), .IN2(n18), .Q(n19) );
  AND2X1 U20 ( .IN1(A[28]), .IN2(n19), .Q(n20) );
  AND2X1 U21 ( .IN1(A[29]), .IN2(n20), .Q(n21) );
  AND2X1 U22 ( .IN1(A[30]), .IN2(n21), .Q(n22) );
  AND2X1 U23 ( .IN1(A[31]), .IN2(n22), .Q(SUM[32]) );
  XOR2X1 U24 ( .IN1(A[31]), .IN2(n22), .Q(SUM[31]) );
  XOR2X1 U25 ( .IN1(A[30]), .IN2(n21), .Q(SUM[30]) );
  XOR2X1 U26 ( .IN1(A[29]), .IN2(n20), .Q(SUM[29]) );
  XOR2X1 U27 ( .IN1(A[28]), .IN2(n19), .Q(SUM[28]) );
  XOR2X1 U28 ( .IN1(A[27]), .IN2(n18), .Q(SUM[27]) );
  XOR2X1 U29 ( .IN1(A[26]), .IN2(n17), .Q(SUM[26]) );
  XOR2X1 U30 ( .IN1(A[25]), .IN2(n16), .Q(SUM[25]) );
  XOR2X1 U31 ( .IN1(A[24]), .IN2(n15), .Q(SUM[24]) );
  XOR2X1 U32 ( .IN1(A[23]), .IN2(n14), .Q(SUM[23]) );
  XOR2X1 U33 ( .IN1(A[22]), .IN2(n13), .Q(SUM[22]) );
  XOR2X1 U34 ( .IN1(A[21]), .IN2(n12), .Q(SUM[21]) );
  XOR2X1 U35 ( .IN1(A[20]), .IN2(n11), .Q(SUM[20]) );
  XOR2X1 U36 ( .IN1(A[19]), .IN2(n10), .Q(SUM[19]) );
  XOR2X1 U37 ( .IN1(A[18]), .IN2(n9), .Q(SUM[18]) );
  XOR2X1 U38 ( .IN1(A[17]), .IN2(n8), .Q(SUM[17]) );
  XOR2X1 U39 ( .IN1(A[16]), .IN2(n7), .Q(SUM[16]) );
  XOR2X1 U40 ( .IN1(A[15]), .IN2(n6), .Q(SUM[15]) );
  XOR2X1 U41 ( .IN1(A[14]), .IN2(n5), .Q(SUM[14]) );
  XOR2X1 U42 ( .IN1(A[13]), .IN2(n4), .Q(SUM[13]) );
  XOR2X1 U43 ( .IN1(A[12]), .IN2(n3), .Q(SUM[12]) );
  XOR2X1 U44 ( .IN1(A[11]), .IN2(n2), .Q(SUM[11]) );
  XOR2X1 U45 ( .IN1(A[10]), .IN2(carry[10]), .Q(SUM[10]) );
  XOR2X1 U46 ( .IN1(A[2]), .IN2(B[2]), .Q(SUM[2]) );
endmodule


module thumb_DW01_add_4 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [32:1] carry;

  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(n2), .CO(carry[4]), .S(SUM[3]) );
  AND2X1 U1 ( .IN1(A[31]), .IN2(n3), .Q(SUM[32]) );
  AND2X1 U2 ( .IN1(A[2]), .IN2(B[2]), .Q(n2) );
  AND2X1 U3 ( .IN1(A[30]), .IN2(n4), .Q(n3) );
  AND2X1 U4 ( .IN1(A[29]), .IN2(n5), .Q(n4) );
  AND2X1 U5 ( .IN1(A[28]), .IN2(n6), .Q(n5) );
  AND2X1 U6 ( .IN1(A[27]), .IN2(n7), .Q(n6) );
  AND2X1 U7 ( .IN1(A[26]), .IN2(n8), .Q(n7) );
  AND2X1 U8 ( .IN1(A[25]), .IN2(n9), .Q(n8) );
  AND2X1 U9 ( .IN1(A[24]), .IN2(n10), .Q(n9) );
  AND2X1 U10 ( .IN1(A[23]), .IN2(n11), .Q(n10) );
  AND2X1 U11 ( .IN1(A[22]), .IN2(n12), .Q(n11) );
  AND2X1 U12 ( .IN1(A[21]), .IN2(n13), .Q(n12) );
  AND2X1 U13 ( .IN1(A[20]), .IN2(n14), .Q(n13) );
  AND2X1 U14 ( .IN1(A[19]), .IN2(n15), .Q(n14) );
  AND2X1 U15 ( .IN1(A[18]), .IN2(n16), .Q(n15) );
  AND2X1 U16 ( .IN1(A[17]), .IN2(n17), .Q(n16) );
  AND2X1 U17 ( .IN1(A[16]), .IN2(n18), .Q(n17) );
  AND2X1 U18 ( .IN1(A[15]), .IN2(n19), .Q(n18) );
  AND2X1 U19 ( .IN1(A[14]), .IN2(n20), .Q(n19) );
  AND2X1 U20 ( .IN1(A[13]), .IN2(n21), .Q(n20) );
  AND2X1 U21 ( .IN1(A[12]), .IN2(n22), .Q(n21) );
  AND2X1 U22 ( .IN1(A[11]), .IN2(n23), .Q(n22) );
  AND2X1 U23 ( .IN1(A[10]), .IN2(carry[10]), .Q(n23) );
  XOR2X1 U24 ( .IN1(A[31]), .IN2(n3), .Q(SUM[31]) );
  XOR2X1 U25 ( .IN1(A[30]), .IN2(n4), .Q(SUM[30]) );
  XOR2X1 U26 ( .IN1(A[29]), .IN2(n5), .Q(SUM[29]) );
  XOR2X1 U27 ( .IN1(A[28]), .IN2(n6), .Q(SUM[28]) );
  XOR2X1 U28 ( .IN1(A[27]), .IN2(n7), .Q(SUM[27]) );
  XOR2X1 U29 ( .IN1(A[26]), .IN2(n8), .Q(SUM[26]) );
  XOR2X1 U30 ( .IN1(A[25]), .IN2(n9), .Q(SUM[25]) );
  XOR2X1 U31 ( .IN1(A[24]), .IN2(n10), .Q(SUM[24]) );
  XOR2X1 U32 ( .IN1(A[23]), .IN2(n11), .Q(SUM[23]) );
  XOR2X1 U33 ( .IN1(A[22]), .IN2(n12), .Q(SUM[22]) );
  XOR2X1 U34 ( .IN1(A[21]), .IN2(n13), .Q(SUM[21]) );
  XOR2X1 U35 ( .IN1(A[20]), .IN2(n14), .Q(SUM[20]) );
  XOR2X1 U36 ( .IN1(A[19]), .IN2(n15), .Q(SUM[19]) );
  XOR2X1 U37 ( .IN1(A[18]), .IN2(n16), .Q(SUM[18]) );
  XOR2X1 U38 ( .IN1(A[17]), .IN2(n17), .Q(SUM[17]) );
  XOR2X1 U39 ( .IN1(A[16]), .IN2(n18), .Q(SUM[16]) );
  XOR2X1 U40 ( .IN1(A[15]), .IN2(n19), .Q(SUM[15]) );
  XOR2X1 U41 ( .IN1(A[14]), .IN2(n20), .Q(SUM[14]) );
  XOR2X1 U42 ( .IN1(A[13]), .IN2(n21), .Q(SUM[13]) );
  XOR2X1 U43 ( .IN1(A[12]), .IN2(n22), .Q(SUM[12]) );
  XOR2X1 U44 ( .IN1(A[11]), .IN2(n23), .Q(SUM[11]) );
  XOR2X1 U45 ( .IN1(A[10]), .IN2(carry[10]), .Q(SUM[10]) );
  XOR2X1 U46 ( .IN1(A[2]), .IN2(B[2]), .Q(SUM[2]) );
endmodule


module thumb_DW01_add_5 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [32:1] carry;

  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(SUM[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module thumb_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29;
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  INVX0 U1 ( .INP(A[1]), .ZN(SUM[1]) );
  XNOR2X1 U2 ( .IN1(A[31]), .IN2(n29), .Q(SUM[31]) );
  NAND2X1 U3 ( .IN1(A[30]), .IN2(n28), .QN(n29) );
  AND2X1 U4 ( .IN1(A[2]), .IN2(A[1]), .Q(n1) );
  AND2X1 U5 ( .IN1(A[3]), .IN2(n1), .Q(n2) );
  AND2X1 U6 ( .IN1(A[4]), .IN2(n2), .Q(n3) );
  AND2X1 U7 ( .IN1(A[5]), .IN2(n3), .Q(n4) );
  AND2X1 U8 ( .IN1(A[6]), .IN2(n4), .Q(n5) );
  AND2X1 U9 ( .IN1(A[7]), .IN2(n5), .Q(n6) );
  AND2X1 U10 ( .IN1(A[8]), .IN2(n6), .Q(n7) );
  AND2X1 U11 ( .IN1(A[9]), .IN2(n7), .Q(n8) );
  AND2X1 U12 ( .IN1(A[10]), .IN2(n8), .Q(n9) );
  AND2X1 U13 ( .IN1(A[11]), .IN2(n9), .Q(n10) );
  AND2X1 U14 ( .IN1(A[12]), .IN2(n10), .Q(n11) );
  AND2X1 U15 ( .IN1(A[13]), .IN2(n11), .Q(n12) );
  AND2X1 U16 ( .IN1(A[14]), .IN2(n12), .Q(n13) );
  AND2X1 U17 ( .IN1(A[15]), .IN2(n13), .Q(n14) );
  AND2X1 U18 ( .IN1(A[16]), .IN2(n14), .Q(n15) );
  AND2X1 U19 ( .IN1(A[17]), .IN2(n15), .Q(n16) );
  AND2X1 U20 ( .IN1(A[18]), .IN2(n16), .Q(n17) );
  AND2X1 U21 ( .IN1(A[19]), .IN2(n17), .Q(n18) );
  AND2X1 U22 ( .IN1(A[20]), .IN2(n18), .Q(n19) );
  AND2X1 U23 ( .IN1(A[21]), .IN2(n19), .Q(n20) );
  AND2X1 U24 ( .IN1(A[22]), .IN2(n20), .Q(n21) );
  AND2X1 U25 ( .IN1(A[23]), .IN2(n21), .Q(n22) );
  AND2X1 U26 ( .IN1(A[24]), .IN2(n22), .Q(n23) );
  AND2X1 U27 ( .IN1(A[25]), .IN2(n23), .Q(n24) );
  AND2X1 U28 ( .IN1(A[26]), .IN2(n24), .Q(n25) );
  AND2X1 U29 ( .IN1(A[27]), .IN2(n25), .Q(n26) );
  AND2X1 U30 ( .IN1(A[28]), .IN2(n26), .Q(n27) );
  AND2X1 U31 ( .IN1(A[29]), .IN2(n27), .Q(n28) );
  XOR2X1 U32 ( .IN1(A[30]), .IN2(n28), .Q(SUM[30]) );
  XOR2X1 U33 ( .IN1(A[29]), .IN2(n27), .Q(SUM[29]) );
  XOR2X1 U34 ( .IN1(A[28]), .IN2(n26), .Q(SUM[28]) );
  XOR2X1 U35 ( .IN1(A[27]), .IN2(n25), .Q(SUM[27]) );
  XOR2X1 U36 ( .IN1(A[26]), .IN2(n24), .Q(SUM[26]) );
  XOR2X1 U37 ( .IN1(A[25]), .IN2(n23), .Q(SUM[25]) );
  XOR2X1 U38 ( .IN1(A[24]), .IN2(n22), .Q(SUM[24]) );
  XOR2X1 U39 ( .IN1(A[23]), .IN2(n21), .Q(SUM[23]) );
  XOR2X1 U40 ( .IN1(A[22]), .IN2(n20), .Q(SUM[22]) );
  XOR2X1 U41 ( .IN1(A[21]), .IN2(n19), .Q(SUM[21]) );
  XOR2X1 U42 ( .IN1(A[20]), .IN2(n18), .Q(SUM[20]) );
  XOR2X1 U43 ( .IN1(A[19]), .IN2(n17), .Q(SUM[19]) );
  XOR2X1 U44 ( .IN1(A[18]), .IN2(n16), .Q(SUM[18]) );
  XOR2X1 U45 ( .IN1(A[17]), .IN2(n15), .Q(SUM[17]) );
  XOR2X1 U46 ( .IN1(A[16]), .IN2(n14), .Q(SUM[16]) );
  XOR2X1 U47 ( .IN1(A[15]), .IN2(n13), .Q(SUM[15]) );
  XOR2X1 U48 ( .IN1(A[14]), .IN2(n12), .Q(SUM[14]) );
  XOR2X1 U49 ( .IN1(A[13]), .IN2(n11), .Q(SUM[13]) );
  XOR2X1 U50 ( .IN1(A[12]), .IN2(n10), .Q(SUM[12]) );
  XOR2X1 U51 ( .IN1(A[11]), .IN2(n9), .Q(SUM[11]) );
  XOR2X1 U52 ( .IN1(A[10]), .IN2(n8), .Q(SUM[10]) );
  XOR2X1 U53 ( .IN1(A[9]), .IN2(n7), .Q(SUM[9]) );
  XOR2X1 U54 ( .IN1(A[8]), .IN2(n6), .Q(SUM[8]) );
  XOR2X1 U55 ( .IN1(A[7]), .IN2(n5), .Q(SUM[7]) );
  XOR2X1 U56 ( .IN1(A[6]), .IN2(n4), .Q(SUM[6]) );
  XOR2X1 U57 ( .IN1(A[5]), .IN2(n3), .Q(SUM[5]) );
  XOR2X1 U58 ( .IN1(A[4]), .IN2(n2), .Q(SUM[4]) );
  XOR2X1 U59 ( .IN1(A[3]), .IN2(n1), .Q(SUM[3]) );
  XOR2X1 U60 ( .IN1(A[2]), .IN2(A[1]), .Q(SUM[2]) );
endmodule


module thumb_DW_leftsh_2 ( A, SH, B );
  input [32:0] A;
  input [7:0] SH;
  output [32:0] B;
  wire   n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n44, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n81, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n118, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n155, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n191, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n306;

  AND2X1 U4 ( .IN1(n41), .IN2(n306), .Q(B[32]) );
  AND2X1 U5 ( .IN1(n40), .IN2(n306), .Q(B[31]) );
  AND2X1 U6 ( .IN1(n39), .IN2(n306), .Q(B[30]) );
  AND2X1 U7 ( .IN1(n38), .IN2(n306), .Q(B[29]) );
  AND2X1 U8 ( .IN1(n37), .IN2(n306), .Q(B[28]) );
  AND2X1 U9 ( .IN1(n36), .IN2(n306), .Q(B[27]) );
  AND2X1 U10 ( .IN1(n35), .IN2(n306), .Q(B[26]) );
  AND2X1 U11 ( .IN1(n34), .IN2(n306), .Q(B[25]) );
  AND2X1 U12 ( .IN1(n33), .IN2(n306), .Q(B[24]) );
  AND2X1 U13 ( .IN1(n32), .IN2(n306), .Q(B[23]) );
  AND2X1 U14 ( .IN1(n31), .IN2(n306), .Q(B[22]) );
  AND2X1 U15 ( .IN1(n30), .IN2(n306), .Q(B[21]) );
  AND2X1 U16 ( .IN1(n29), .IN2(n306), .Q(B[20]) );
  AND2X1 U17 ( .IN1(n28), .IN2(n306), .Q(B[19]) );
  AND2X1 U18 ( .IN1(n27), .IN2(n306), .Q(B[18]) );
  AND2X1 U19 ( .IN1(n26), .IN2(n306), .Q(B[17]) );
  AND2X1 U20 ( .IN1(n25), .IN2(n306), .Q(B[16]) );
  AND2X1 U21 ( .IN1(n24), .IN2(n306), .Q(B[15]) );
  AND2X1 U22 ( .IN1(n23), .IN2(n306), .Q(B[14]) );
  AND2X1 U23 ( .IN1(n22), .IN2(n306), .Q(B[13]) );
  AND2X1 U24 ( .IN1(n21), .IN2(n306), .Q(B[12]) );
  AND2X1 U25 ( .IN1(n20), .IN2(n306), .Q(B[11]) );
  AND2X1 U26 ( .IN1(n19), .IN2(n306), .Q(B[10]) );
  AND2X1 U27 ( .IN1(n18), .IN2(n306), .Q(B[9]) );
  AND2X1 U28 ( .IN1(n17), .IN2(n306), .Q(B[8]) );
  AND2X1 U29 ( .IN1(n16), .IN2(n306), .Q(B[7]) );
  AND2X1 U30 ( .IN1(n15), .IN2(n306), .Q(B[6]) );
  AND2X1 U31 ( .IN1(n14), .IN2(n306), .Q(B[5]) );
  AND2X1 U32 ( .IN1(n13), .IN2(n306), .Q(B[4]) );
  AND2X1 U33 ( .IN1(n12), .IN2(n306), .Q(B[3]) );
  AND2X1 U34 ( .IN1(n11), .IN2(n306), .Q(B[2]) );
  AND2X1 U35 ( .IN1(n10), .IN2(n306), .Q(B[1]) );
  AND2X1 U36 ( .IN1(n9), .IN2(n306), .Q(B[0]) );
  AO22X1 U41 ( .IN1(SH[5]), .IN2(n46), .IN3(n78), .IN4(n7), .Q(n41) );
  AND2X1 U42 ( .IN1(n77), .IN2(n7), .Q(n40) );
  AND2X1 U43 ( .IN1(n76), .IN2(n7), .Q(n39) );
  AND2X1 U44 ( .IN1(n75), .IN2(n7), .Q(n38) );
  AND2X1 U45 ( .IN1(n74), .IN2(n7), .Q(n37) );
  AND2X1 U46 ( .IN1(n73), .IN2(n7), .Q(n36) );
  AND2X1 U47 ( .IN1(n72), .IN2(n7), .Q(n35) );
  AND2X1 U48 ( .IN1(n71), .IN2(n7), .Q(n34) );
  AND2X1 U49 ( .IN1(n70), .IN2(n7), .Q(n33) );
  AND2X1 U50 ( .IN1(n69), .IN2(n7), .Q(n32) );
  AND2X1 U51 ( .IN1(n68), .IN2(n7), .Q(n31) );
  AND2X1 U52 ( .IN1(n67), .IN2(n7), .Q(n30) );
  AND2X1 U53 ( .IN1(n66), .IN2(n7), .Q(n29) );
  AND2X1 U54 ( .IN1(n65), .IN2(n7), .Q(n28) );
  AND2X1 U55 ( .IN1(n64), .IN2(n7), .Q(n27) );
  AND2X1 U56 ( .IN1(n63), .IN2(n7), .Q(n26) );
  AND2X1 U57 ( .IN1(n62), .IN2(n7), .Q(n25) );
  AND2X1 U58 ( .IN1(n61), .IN2(n7), .Q(n24) );
  AND2X1 U59 ( .IN1(n60), .IN2(n7), .Q(n23) );
  AND2X1 U60 ( .IN1(n59), .IN2(n7), .Q(n22) );
  AND2X1 U61 ( .IN1(n58), .IN2(n7), .Q(n21) );
  AND2X1 U62 ( .IN1(n57), .IN2(n7), .Q(n20) );
  AND2X1 U63 ( .IN1(n56), .IN2(n7), .Q(n19) );
  AND2X1 U64 ( .IN1(n55), .IN2(n7), .Q(n18) );
  AND2X1 U65 ( .IN1(n54), .IN2(n7), .Q(n17) );
  AND2X1 U66 ( .IN1(n53), .IN2(n7), .Q(n16) );
  AND2X1 U67 ( .IN1(n52), .IN2(n7), .Q(n15) );
  AND2X1 U68 ( .IN1(n51), .IN2(n7), .Q(n14) );
  AND2X1 U69 ( .IN1(n50), .IN2(n7), .Q(n13) );
  AND2X1 U70 ( .IN1(n49), .IN2(n7), .Q(n12) );
  AND2X1 U71 ( .IN1(n48), .IN2(n7), .Q(n11) );
  AND2X1 U72 ( .IN1(n47), .IN2(n7), .Q(n10) );
  AND2X1 U73 ( .IN1(n46), .IN2(n7), .Q(n9) );
  AO22X1 U78 ( .IN1(n44), .IN2(n115), .IN3(n99), .IN4(SH[4]), .Q(n78) );
  AO22X1 U79 ( .IN1(SH[4]), .IN2(n98), .IN3(n114), .IN4(n44), .Q(n77) );
  AO22X1 U80 ( .IN1(SH[4]), .IN2(n97), .IN3(n113), .IN4(n44), .Q(n76) );
  AO22X1 U81 ( .IN1(SH[4]), .IN2(n96), .IN3(n112), .IN4(n44), .Q(n75) );
  AO22X1 U82 ( .IN1(SH[4]), .IN2(n95), .IN3(n111), .IN4(n44), .Q(n74) );
  AO22X1 U83 ( .IN1(SH[4]), .IN2(n94), .IN3(n110), .IN4(n44), .Q(n73) );
  AO22X1 U84 ( .IN1(SH[4]), .IN2(n93), .IN3(n109), .IN4(n44), .Q(n72) );
  AO22X1 U85 ( .IN1(SH[4]), .IN2(n92), .IN3(n108), .IN4(n44), .Q(n71) );
  AO22X1 U86 ( .IN1(SH[4]), .IN2(n91), .IN3(n107), .IN4(n44), .Q(n70) );
  AO22X1 U87 ( .IN1(SH[4]), .IN2(n90), .IN3(n106), .IN4(n44), .Q(n69) );
  AO22X1 U88 ( .IN1(SH[4]), .IN2(n89), .IN3(n105), .IN4(n44), .Q(n68) );
  AO22X1 U89 ( .IN1(SH[4]), .IN2(n88), .IN3(n104), .IN4(n44), .Q(n67) );
  AO22X1 U90 ( .IN1(SH[4]), .IN2(n87), .IN3(n103), .IN4(n44), .Q(n66) );
  AO22X1 U91 ( .IN1(SH[4]), .IN2(n86), .IN3(n102), .IN4(n44), .Q(n65) );
  AO22X1 U92 ( .IN1(SH[4]), .IN2(n85), .IN3(n101), .IN4(n44), .Q(n64) );
  AO22X1 U93 ( .IN1(SH[4]), .IN2(n84), .IN3(n100), .IN4(n44), .Q(n63) );
  AO22X1 U94 ( .IN1(SH[4]), .IN2(n83), .IN3(n99), .IN4(n44), .Q(n62) );
  AND2X1 U95 ( .IN1(n98), .IN2(n44), .Q(n61) );
  AND2X1 U96 ( .IN1(n97), .IN2(n44), .Q(n60) );
  AND2X1 U97 ( .IN1(n96), .IN2(n44), .Q(n59) );
  AND2X1 U98 ( .IN1(n95), .IN2(n44), .Q(n58) );
  AND2X1 U99 ( .IN1(n94), .IN2(n44), .Q(n57) );
  AND2X1 U100 ( .IN1(n93), .IN2(n44), .Q(n56) );
  AND2X1 U101 ( .IN1(n92), .IN2(n44), .Q(n55) );
  AND2X1 U102 ( .IN1(n91), .IN2(n44), .Q(n54) );
  AND2X1 U103 ( .IN1(n90), .IN2(n44), .Q(n53) );
  AND2X1 U104 ( .IN1(n89), .IN2(n44), .Q(n52) );
  AND2X1 U105 ( .IN1(n88), .IN2(n44), .Q(n51) );
  AND2X1 U106 ( .IN1(n87), .IN2(n44), .Q(n50) );
  AND2X1 U107 ( .IN1(n86), .IN2(n44), .Q(n49) );
  AND2X1 U108 ( .IN1(n85), .IN2(n44), .Q(n48) );
  AND2X1 U109 ( .IN1(n84), .IN2(n44), .Q(n47) );
  AND2X1 U110 ( .IN1(n83), .IN2(n44), .Q(n46) );
  AO22X1 U115 ( .IN1(n81), .IN2(n152), .IN3(n144), .IN4(SH[3]), .Q(n115) );
  AO22X1 U116 ( .IN1(SH[3]), .IN2(n143), .IN3(n151), .IN4(n81), .Q(n114) );
  AO22X1 U117 ( .IN1(SH[3]), .IN2(n142), .IN3(n150), .IN4(n81), .Q(n113) );
  AO22X1 U118 ( .IN1(SH[3]), .IN2(n141), .IN3(n149), .IN4(n81), .Q(n112) );
  AO22X1 U119 ( .IN1(SH[3]), .IN2(n140), .IN3(n148), .IN4(n81), .Q(n111) );
  AO22X1 U120 ( .IN1(SH[3]), .IN2(n139), .IN3(n147), .IN4(n81), .Q(n110) );
  AO22X1 U121 ( .IN1(SH[3]), .IN2(n138), .IN3(n146), .IN4(n81), .Q(n109) );
  AO22X1 U122 ( .IN1(SH[3]), .IN2(n137), .IN3(n145), .IN4(n81), .Q(n108) );
  AO22X1 U123 ( .IN1(SH[3]), .IN2(n136), .IN3(n144), .IN4(n81), .Q(n107) );
  AO22X1 U124 ( .IN1(SH[3]), .IN2(n135), .IN3(n143), .IN4(n81), .Q(n106) );
  AO22X1 U125 ( .IN1(SH[3]), .IN2(n134), .IN3(n142), .IN4(n81), .Q(n105) );
  AO22X1 U126 ( .IN1(SH[3]), .IN2(n133), .IN3(n141), .IN4(n81), .Q(n104) );
  AO22X1 U127 ( .IN1(SH[3]), .IN2(n132), .IN3(n140), .IN4(n81), .Q(n103) );
  AO22X1 U128 ( .IN1(SH[3]), .IN2(n131), .IN3(n139), .IN4(n81), .Q(n102) );
  AO22X1 U129 ( .IN1(SH[3]), .IN2(n130), .IN3(n138), .IN4(n81), .Q(n101) );
  AO22X1 U130 ( .IN1(SH[3]), .IN2(n129), .IN3(n137), .IN4(n81), .Q(n100) );
  AO22X1 U131 ( .IN1(SH[3]), .IN2(n128), .IN3(n136), .IN4(n81), .Q(n99) );
  AO22X1 U132 ( .IN1(SH[3]), .IN2(n127), .IN3(n135), .IN4(n81), .Q(n98) );
  AO22X1 U133 ( .IN1(SH[3]), .IN2(n126), .IN3(n134), .IN4(n81), .Q(n97) );
  AO22X1 U134 ( .IN1(SH[3]), .IN2(n125), .IN3(n133), .IN4(n81), .Q(n96) );
  AO22X1 U135 ( .IN1(SH[3]), .IN2(n124), .IN3(n132), .IN4(n81), .Q(n95) );
  AO22X1 U136 ( .IN1(SH[3]), .IN2(n123), .IN3(n131), .IN4(n81), .Q(n94) );
  AO22X1 U137 ( .IN1(SH[3]), .IN2(n122), .IN3(n130), .IN4(n81), .Q(n93) );
  AO22X1 U138 ( .IN1(SH[3]), .IN2(n121), .IN3(n129), .IN4(n81), .Q(n92) );
  AO22X1 U139 ( .IN1(SH[3]), .IN2(n120), .IN3(n128), .IN4(n81), .Q(n91) );
  AND2X1 U140 ( .IN1(n127), .IN2(n81), .Q(n90) );
  AND2X1 U141 ( .IN1(n126), .IN2(n81), .Q(n89) );
  AND2X1 U142 ( .IN1(n125), .IN2(n81), .Q(n88) );
  AND2X1 U143 ( .IN1(n124), .IN2(n81), .Q(n87) );
  AND2X1 U144 ( .IN1(n123), .IN2(n81), .Q(n86) );
  AND2X1 U145 ( .IN1(n122), .IN2(n81), .Q(n85) );
  AND2X1 U146 ( .IN1(n121), .IN2(n81), .Q(n84) );
  AND2X1 U147 ( .IN1(n120), .IN2(n81), .Q(n83) );
  AO22X1 U152 ( .IN1(n118), .IN2(n189), .IN3(n185), .IN4(SH[2]), .Q(n152) );
  AO22X1 U153 ( .IN1(SH[2]), .IN2(n184), .IN3(n188), .IN4(n118), .Q(n151) );
  AO22X1 U154 ( .IN1(SH[2]), .IN2(n183), .IN3(n187), .IN4(n118), .Q(n150) );
  AO22X1 U155 ( .IN1(SH[2]), .IN2(n182), .IN3(n186), .IN4(n118), .Q(n149) );
  AO22X1 U156 ( .IN1(SH[2]), .IN2(n181), .IN3(n185), .IN4(n118), .Q(n148) );
  AO22X1 U157 ( .IN1(SH[2]), .IN2(n180), .IN3(n184), .IN4(n118), .Q(n147) );
  AO22X1 U158 ( .IN1(SH[2]), .IN2(n179), .IN3(n183), .IN4(n118), .Q(n146) );
  AO22X1 U159 ( .IN1(SH[2]), .IN2(n178), .IN3(n182), .IN4(n118), .Q(n145) );
  AO22X1 U160 ( .IN1(SH[2]), .IN2(n177), .IN3(n181), .IN4(n118), .Q(n144) );
  AO22X1 U161 ( .IN1(SH[2]), .IN2(n176), .IN3(n180), .IN4(n118), .Q(n143) );
  AO22X1 U162 ( .IN1(SH[2]), .IN2(n175), .IN3(n179), .IN4(n118), .Q(n142) );
  AO22X1 U163 ( .IN1(SH[2]), .IN2(n174), .IN3(n178), .IN4(n118), .Q(n141) );
  AO22X1 U164 ( .IN1(SH[2]), .IN2(n173), .IN3(n177), .IN4(n118), .Q(n140) );
  AO22X1 U165 ( .IN1(SH[2]), .IN2(n172), .IN3(n176), .IN4(n118), .Q(n139) );
  AO22X1 U166 ( .IN1(SH[2]), .IN2(n171), .IN3(n175), .IN4(n118), .Q(n138) );
  AO22X1 U167 ( .IN1(SH[2]), .IN2(n170), .IN3(n174), .IN4(n118), .Q(n137) );
  AO22X1 U168 ( .IN1(SH[2]), .IN2(n169), .IN3(n173), .IN4(n118), .Q(n136) );
  AO22X1 U169 ( .IN1(SH[2]), .IN2(n168), .IN3(n172), .IN4(n118), .Q(n135) );
  AO22X1 U170 ( .IN1(SH[2]), .IN2(n167), .IN3(n171), .IN4(n118), .Q(n134) );
  AO22X1 U171 ( .IN1(SH[2]), .IN2(n166), .IN3(n170), .IN4(n118), .Q(n133) );
  AO22X1 U172 ( .IN1(SH[2]), .IN2(n165), .IN3(n169), .IN4(n118), .Q(n132) );
  AO22X1 U173 ( .IN1(SH[2]), .IN2(n164), .IN3(n168), .IN4(n118), .Q(n131) );
  AO22X1 U174 ( .IN1(SH[2]), .IN2(n163), .IN3(n167), .IN4(n118), .Q(n130) );
  AO22X1 U175 ( .IN1(SH[2]), .IN2(n162), .IN3(n166), .IN4(n118), .Q(n129) );
  AO22X1 U176 ( .IN1(SH[2]), .IN2(n161), .IN3(n165), .IN4(n118), .Q(n128) );
  AO22X1 U177 ( .IN1(SH[2]), .IN2(n160), .IN3(n164), .IN4(n118), .Q(n127) );
  AO22X1 U178 ( .IN1(SH[2]), .IN2(n159), .IN3(n163), .IN4(n118), .Q(n126) );
  AO22X1 U179 ( .IN1(SH[2]), .IN2(n158), .IN3(n162), .IN4(n118), .Q(n125) );
  AO22X1 U180 ( .IN1(SH[2]), .IN2(n157), .IN3(n161), .IN4(n118), .Q(n124) );
  AND2X1 U181 ( .IN1(n160), .IN2(n118), .Q(n123) );
  AND2X1 U182 ( .IN1(n159), .IN2(n118), .Q(n122) );
  AND2X1 U183 ( .IN1(n158), .IN2(n118), .Q(n121) );
  AND2X1 U184 ( .IN1(n157), .IN2(n118), .Q(n120) );
  AO22X1 U189 ( .IN1(n225), .IN2(n155), .IN3(n223), .IN4(SH[1]), .Q(n189) );
  AO22X1 U190 ( .IN1(SH[1]), .IN2(n222), .IN3(n224), .IN4(n155), .Q(n188) );
  AO22X1 U191 ( .IN1(SH[1]), .IN2(n221), .IN3(n223), .IN4(n155), .Q(n187) );
  AO22X1 U192 ( .IN1(SH[1]), .IN2(n220), .IN3(n222), .IN4(n155), .Q(n186) );
  AO22X1 U193 ( .IN1(SH[1]), .IN2(n219), .IN3(n221), .IN4(n155), .Q(n185) );
  AO22X1 U194 ( .IN1(SH[1]), .IN2(n218), .IN3(n220), .IN4(n155), .Q(n184) );
  AO22X1 U195 ( .IN1(SH[1]), .IN2(n217), .IN3(n219), .IN4(n155), .Q(n183) );
  AO22X1 U196 ( .IN1(SH[1]), .IN2(n216), .IN3(n218), .IN4(n155), .Q(n182) );
  AO22X1 U197 ( .IN1(SH[1]), .IN2(n215), .IN3(n217), .IN4(n155), .Q(n181) );
  AO22X1 U198 ( .IN1(SH[1]), .IN2(n214), .IN3(n216), .IN4(n155), .Q(n180) );
  AO22X1 U199 ( .IN1(SH[1]), .IN2(n213), .IN3(n215), .IN4(n155), .Q(n179) );
  AO22X1 U200 ( .IN1(SH[1]), .IN2(n212), .IN3(n214), .IN4(n155), .Q(n178) );
  AO22X1 U201 ( .IN1(SH[1]), .IN2(n211), .IN3(n213), .IN4(n155), .Q(n177) );
  AO22X1 U202 ( .IN1(SH[1]), .IN2(n210), .IN3(n212), .IN4(n155), .Q(n176) );
  AO22X1 U203 ( .IN1(SH[1]), .IN2(n209), .IN3(n211), .IN4(n155), .Q(n175) );
  AO22X1 U204 ( .IN1(SH[1]), .IN2(n208), .IN3(n210), .IN4(n155), .Q(n174) );
  AO22X1 U205 ( .IN1(SH[1]), .IN2(n207), .IN3(n209), .IN4(n155), .Q(n173) );
  AO22X1 U206 ( .IN1(SH[1]), .IN2(n206), .IN3(n208), .IN4(n155), .Q(n172) );
  AO22X1 U207 ( .IN1(SH[1]), .IN2(n205), .IN3(n207), .IN4(n155), .Q(n171) );
  AO22X1 U208 ( .IN1(SH[1]), .IN2(n204), .IN3(n206), .IN4(n155), .Q(n170) );
  AO22X1 U209 ( .IN1(SH[1]), .IN2(n203), .IN3(n205), .IN4(n155), .Q(n169) );
  AO22X1 U210 ( .IN1(SH[1]), .IN2(n202), .IN3(n204), .IN4(n155), .Q(n168) );
  AO22X1 U211 ( .IN1(SH[1]), .IN2(n201), .IN3(n203), .IN4(n155), .Q(n167) );
  AO22X1 U212 ( .IN1(SH[1]), .IN2(n200), .IN3(n202), .IN4(n155), .Q(n166) );
  AO22X1 U213 ( .IN1(SH[1]), .IN2(n199), .IN3(n201), .IN4(n155), .Q(n165) );
  AO22X1 U214 ( .IN1(SH[1]), .IN2(n198), .IN3(n200), .IN4(n155), .Q(n164) );
  AO22X1 U215 ( .IN1(SH[1]), .IN2(n197), .IN3(n199), .IN4(n155), .Q(n163) );
  AO22X1 U216 ( .IN1(SH[1]), .IN2(n196), .IN3(n198), .IN4(n155), .Q(n162) );
  AO22X1 U217 ( .IN1(SH[1]), .IN2(n195), .IN3(n197), .IN4(n155), .Q(n161) );
  AO22X1 U218 ( .IN1(SH[1]), .IN2(n194), .IN3(n196), .IN4(n155), .Q(n160) );
  AO22X1 U219 ( .IN1(SH[1]), .IN2(n193), .IN3(n195), .IN4(n155), .Q(n159) );
  AND2X1 U220 ( .IN1(n194), .IN2(n155), .Q(n158) );
  AND2X1 U221 ( .IN1(n193), .IN2(n155), .Q(n157) );
  AND2X1 U225 ( .IN1(SH[0]), .IN2(A[31]), .Q(n225) );
  AO22X1 U226 ( .IN1(A[30]), .IN2(SH[0]), .IN3(n191), .IN4(A[31]), .Q(n224) );
  AO22X1 U227 ( .IN1(A[29]), .IN2(SH[0]), .IN3(n191), .IN4(A[30]), .Q(n223) );
  AO22X1 U228 ( .IN1(A[28]), .IN2(SH[0]), .IN3(n191), .IN4(A[29]), .Q(n222) );
  AO22X1 U229 ( .IN1(A[27]), .IN2(SH[0]), .IN3(n191), .IN4(A[28]), .Q(n221) );
  AO22X1 U230 ( .IN1(A[26]), .IN2(SH[0]), .IN3(n191), .IN4(A[27]), .Q(n220) );
  AO22X1 U231 ( .IN1(A[25]), .IN2(SH[0]), .IN3(n191), .IN4(A[26]), .Q(n219) );
  AO22X1 U232 ( .IN1(A[24]), .IN2(SH[0]), .IN3(n191), .IN4(A[25]), .Q(n218) );
  AO22X1 U233 ( .IN1(A[23]), .IN2(SH[0]), .IN3(n191), .IN4(A[24]), .Q(n217) );
  AO22X1 U234 ( .IN1(A[22]), .IN2(SH[0]), .IN3(n191), .IN4(A[23]), .Q(n216) );
  AO22X1 U235 ( .IN1(A[21]), .IN2(SH[0]), .IN3(n191), .IN4(A[22]), .Q(n215) );
  AO22X1 U236 ( .IN1(A[20]), .IN2(SH[0]), .IN3(n191), .IN4(A[21]), .Q(n214) );
  AO22X1 U237 ( .IN1(A[19]), .IN2(SH[0]), .IN3(n191), .IN4(A[20]), .Q(n213) );
  AO22X1 U238 ( .IN1(A[18]), .IN2(SH[0]), .IN3(n191), .IN4(A[19]), .Q(n212) );
  AO22X1 U239 ( .IN1(A[17]), .IN2(SH[0]), .IN3(n191), .IN4(A[18]), .Q(n211) );
  AO22X1 U240 ( .IN1(A[16]), .IN2(SH[0]), .IN3(n191), .IN4(A[17]), .Q(n210) );
  AO22X1 U241 ( .IN1(A[15]), .IN2(SH[0]), .IN3(n191), .IN4(A[16]), .Q(n209) );
  AO22X1 U242 ( .IN1(A[14]), .IN2(SH[0]), .IN3(n191), .IN4(A[15]), .Q(n208) );
  AO22X1 U243 ( .IN1(A[13]), .IN2(SH[0]), .IN3(n191), .IN4(A[14]), .Q(n207) );
  AO22X1 U244 ( .IN1(A[12]), .IN2(SH[0]), .IN3(n191), .IN4(A[13]), .Q(n206) );
  AO22X1 U245 ( .IN1(A[11]), .IN2(SH[0]), .IN3(n191), .IN4(A[12]), .Q(n205) );
  AO22X1 U246 ( .IN1(A[10]), .IN2(SH[0]), .IN3(n191), .IN4(A[11]), .Q(n204) );
  AO22X1 U247 ( .IN1(A[9]), .IN2(SH[0]), .IN3(n191), .IN4(A[10]), .Q(n203) );
  AO22X1 U248 ( .IN1(A[8]), .IN2(SH[0]), .IN3(n191), .IN4(A[9]), .Q(n202) );
  AO22X1 U249 ( .IN1(A[7]), .IN2(SH[0]), .IN3(n191), .IN4(A[8]), .Q(n201) );
  AO22X1 U250 ( .IN1(A[6]), .IN2(SH[0]), .IN3(n191), .IN4(A[7]), .Q(n200) );
  AO22X1 U251 ( .IN1(A[5]), .IN2(SH[0]), .IN3(n191), .IN4(A[6]), .Q(n199) );
  AO22X1 U252 ( .IN1(A[4]), .IN2(SH[0]), .IN3(n191), .IN4(A[5]), .Q(n198) );
  AO22X1 U253 ( .IN1(A[3]), .IN2(SH[0]), .IN3(n191), .IN4(A[4]), .Q(n197) );
  AO22X1 U254 ( .IN1(A[2]), .IN2(SH[0]), .IN3(n191), .IN4(A[3]), .Q(n196) );
  AO22X1 U255 ( .IN1(A[1]), .IN2(SH[0]), .IN3(n191), .IN4(A[2]), .Q(n195) );
  AO22X1 U256 ( .IN1(A[0]), .IN2(SH[0]), .IN3(n191), .IN4(A[1]), .Q(n194) );
  AND2X1 U257 ( .IN1(n191), .IN2(A[0]), .Q(n193) );
  INVX0 U263 ( .INP(SH[1]), .ZN(n155) );
  INVX0 U264 ( .INP(SH[0]), .ZN(n191) );
  INVX0 U265 ( .INP(SH[2]), .ZN(n118) );
  INVX0 U266 ( .INP(SH[3]), .ZN(n81) );
  INVX0 U267 ( .INP(SH[4]), .ZN(n44) );
  INVX0 U268 ( .INP(SH[5]), .ZN(n7) );
  NOR2X0 U269 ( .IN1(SH[7]), .IN2(SH[6]), .QN(n306) );
endmodule


module thumb_DW_rightsh_3 ( A, DATA_TC, SH, B );
  input [32:0] A;
  input [4:0] SH;
  output [32:0] B;
  input DATA_TC;
  wire   n1, n17, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163;

  MUX21X1 U33 ( .IN1(n41), .IN2(n57), .S(SH[4]), .Q(B[16]) );
  MUX21X1 U34 ( .IN1(n40), .IN2(n56), .S(SH[4]), .Q(B[15]) );
  MUX21X1 U35 ( .IN1(n39), .IN2(n55), .S(SH[4]), .Q(B[14]) );
  MUX21X1 U36 ( .IN1(n38), .IN2(n54), .S(SH[4]), .Q(B[13]) );
  MUX21X1 U37 ( .IN1(n37), .IN2(n53), .S(SH[4]), .Q(B[12]) );
  MUX21X1 U38 ( .IN1(n36), .IN2(n52), .S(SH[4]), .Q(B[11]) );
  MUX21X1 U39 ( .IN1(n35), .IN2(n51), .S(SH[4]), .Q(B[10]) );
  MUX21X1 U40 ( .IN1(n34), .IN2(n50), .S(SH[4]), .Q(B[9]) );
  MUX21X1 U41 ( .IN1(n33), .IN2(n49), .S(SH[4]), .Q(B[8]) );
  MUX21X1 U42 ( .IN1(n32), .IN2(n48), .S(SH[4]), .Q(B[7]) );
  MUX21X1 U43 ( .IN1(n31), .IN2(n47), .S(SH[4]), .Q(B[6]) );
  MUX21X1 U44 ( .IN1(n30), .IN2(n46), .S(SH[4]), .Q(B[5]) );
  MUX21X1 U45 ( .IN1(n29), .IN2(n45), .S(SH[4]), .Q(B[4]) );
  MUX21X1 U46 ( .IN1(n28), .IN2(n44), .S(SH[4]), .Q(B[3]) );
  MUX21X1 U47 ( .IN1(n27), .IN2(n43), .S(SH[4]), .Q(B[2]) );
  MUX21X1 U48 ( .IN1(n26), .IN2(n42), .S(SH[4]), .Q(B[1]) );
  MUX21X1 U49 ( .IN1(n25), .IN2(n41), .S(SH[4]), .Q(B[0]) );
  MUX21X1 U66 ( .IN1(n86), .IN2(n94), .S(SH[3]), .Q(n49) );
  MUX21X1 U67 ( .IN1(n85), .IN2(n93), .S(SH[3]), .Q(n48) );
  MUX21X1 U68 ( .IN1(n84), .IN2(n92), .S(SH[3]), .Q(n47) );
  MUX21X1 U69 ( .IN1(n83), .IN2(n91), .S(SH[3]), .Q(n46) );
  MUX21X1 U70 ( .IN1(n82), .IN2(n90), .S(SH[3]), .Q(n45) );
  MUX21X1 U71 ( .IN1(n81), .IN2(n89), .S(SH[3]), .Q(n44) );
  MUX21X1 U72 ( .IN1(n80), .IN2(n88), .S(SH[3]), .Q(n43) );
  MUX21X1 U73 ( .IN1(n79), .IN2(n87), .S(SH[3]), .Q(n42) );
  MUX21X1 U74 ( .IN1(n78), .IN2(n86), .S(SH[3]), .Q(n41) );
  MUX21X1 U75 ( .IN1(n77), .IN2(n85), .S(SH[3]), .Q(n40) );
  MUX21X1 U76 ( .IN1(n76), .IN2(n84), .S(SH[3]), .Q(n39) );
  MUX21X1 U77 ( .IN1(n75), .IN2(n83), .S(SH[3]), .Q(n38) );
  MUX21X1 U78 ( .IN1(n74), .IN2(n82), .S(SH[3]), .Q(n37) );
  MUX21X1 U79 ( .IN1(n73), .IN2(n81), .S(SH[3]), .Q(n36) );
  MUX21X1 U80 ( .IN1(n72), .IN2(n80), .S(SH[3]), .Q(n35) );
  MUX21X1 U81 ( .IN1(n71), .IN2(n79), .S(SH[3]), .Q(n34) );
  MUX21X1 U82 ( .IN1(n70), .IN2(n78), .S(SH[3]), .Q(n33) );
  MUX21X1 U83 ( .IN1(n69), .IN2(n77), .S(SH[3]), .Q(n32) );
  MUX21X1 U84 ( .IN1(n68), .IN2(n76), .S(SH[3]), .Q(n31) );
  MUX21X1 U85 ( .IN1(n67), .IN2(n75), .S(SH[3]), .Q(n30) );
  MUX21X1 U86 ( .IN1(n66), .IN2(n74), .S(SH[3]), .Q(n29) );
  MUX21X1 U87 ( .IN1(n65), .IN2(n73), .S(SH[3]), .Q(n28) );
  MUX21X1 U88 ( .IN1(n64), .IN2(n72), .S(SH[3]), .Q(n27) );
  MUX21X1 U89 ( .IN1(n63), .IN2(n71), .S(SH[3]), .Q(n26) );
  MUX21X1 U90 ( .IN1(n62), .IN2(n70), .S(SH[3]), .Q(n25) );
  MUX21X1 U99 ( .IN1(n125), .IN2(n129), .S(SH[2]), .Q(n90) );
  MUX21X1 U100 ( .IN1(n124), .IN2(n128), .S(SH[2]), .Q(n89) );
  MUX21X1 U101 ( .IN1(n123), .IN2(n127), .S(SH[2]), .Q(n88) );
  MUX21X1 U102 ( .IN1(n122), .IN2(n126), .S(SH[2]), .Q(n87) );
  MUX21X1 U103 ( .IN1(n121), .IN2(n125), .S(SH[2]), .Q(n86) );
  MUX21X1 U104 ( .IN1(n120), .IN2(n124), .S(SH[2]), .Q(n85) );
  MUX21X1 U105 ( .IN1(n119), .IN2(n123), .S(SH[2]), .Q(n84) );
  MUX21X1 U106 ( .IN1(n118), .IN2(n122), .S(SH[2]), .Q(n83) );
  MUX21X1 U107 ( .IN1(n117), .IN2(n121), .S(SH[2]), .Q(n82) );
  MUX21X1 U108 ( .IN1(n116), .IN2(n120), .S(SH[2]), .Q(n81) );
  MUX21X1 U109 ( .IN1(n115), .IN2(n119), .S(SH[2]), .Q(n80) );
  MUX21X1 U110 ( .IN1(n114), .IN2(n118), .S(SH[2]), .Q(n79) );
  MUX21X1 U111 ( .IN1(n113), .IN2(n117), .S(SH[2]), .Q(n78) );
  MUX21X1 U112 ( .IN1(n112), .IN2(n116), .S(SH[2]), .Q(n77) );
  MUX21X1 U113 ( .IN1(n111), .IN2(n115), .S(SH[2]), .Q(n76) );
  MUX21X1 U114 ( .IN1(n110), .IN2(n114), .S(SH[2]), .Q(n75) );
  MUX21X1 U115 ( .IN1(n109), .IN2(n113), .S(SH[2]), .Q(n74) );
  MUX21X1 U116 ( .IN1(n108), .IN2(n112), .S(SH[2]), .Q(n73) );
  MUX21X1 U117 ( .IN1(n107), .IN2(n111), .S(SH[2]), .Q(n72) );
  MUX21X1 U118 ( .IN1(n106), .IN2(n110), .S(SH[2]), .Q(n71) );
  MUX21X1 U119 ( .IN1(n105), .IN2(n109), .S(SH[2]), .Q(n70) );
  MUX21X1 U120 ( .IN1(n104), .IN2(n108), .S(SH[2]), .Q(n69) );
  MUX21X1 U121 ( .IN1(n103), .IN2(n107), .S(SH[2]), .Q(n68) );
  MUX21X1 U122 ( .IN1(n102), .IN2(n106), .S(SH[2]), .Q(n67) );
  MUX21X1 U123 ( .IN1(n101), .IN2(n105), .S(SH[2]), .Q(n66) );
  MUX21X1 U124 ( .IN1(n100), .IN2(n104), .S(SH[2]), .Q(n65) );
  MUX21X1 U125 ( .IN1(n99), .IN2(n103), .S(SH[2]), .Q(n64) );
  MUX21X1 U126 ( .IN1(n98), .IN2(n102), .S(SH[2]), .Q(n63) );
  MUX21X1 U127 ( .IN1(n97), .IN2(n101), .S(SH[2]), .Q(n62) );
  MUX21X1 U132 ( .IN1(n161), .IN2(n163), .S(SH[1]), .Q(n127) );
  MUX21X1 U133 ( .IN1(n160), .IN2(n162), .S(SH[1]), .Q(n126) );
  MUX21X1 U134 ( .IN1(n159), .IN2(n161), .S(SH[1]), .Q(n125) );
  MUX21X1 U135 ( .IN1(n158), .IN2(n160), .S(SH[1]), .Q(n124) );
  MUX21X1 U136 ( .IN1(n157), .IN2(n159), .S(SH[1]), .Q(n123) );
  MUX21X1 U137 ( .IN1(n156), .IN2(n158), .S(SH[1]), .Q(n122) );
  MUX21X1 U138 ( .IN1(n155), .IN2(n157), .S(SH[1]), .Q(n121) );
  MUX21X1 U139 ( .IN1(n154), .IN2(n156), .S(SH[1]), .Q(n120) );
  MUX21X1 U140 ( .IN1(n153), .IN2(n155), .S(SH[1]), .Q(n119) );
  MUX21X1 U141 ( .IN1(n152), .IN2(n154), .S(SH[1]), .Q(n118) );
  MUX21X1 U142 ( .IN1(n151), .IN2(n153), .S(SH[1]), .Q(n117) );
  MUX21X1 U143 ( .IN1(n150), .IN2(n152), .S(SH[1]), .Q(n116) );
  MUX21X1 U144 ( .IN1(n149), .IN2(n151), .S(SH[1]), .Q(n115) );
  MUX21X1 U145 ( .IN1(n148), .IN2(n150), .S(SH[1]), .Q(n114) );
  MUX21X1 U146 ( .IN1(n147), .IN2(n149), .S(SH[1]), .Q(n113) );
  MUX21X1 U147 ( .IN1(n146), .IN2(n148), .S(SH[1]), .Q(n112) );
  MUX21X1 U148 ( .IN1(n145), .IN2(n147), .S(SH[1]), .Q(n111) );
  MUX21X1 U149 ( .IN1(n144), .IN2(n146), .S(SH[1]), .Q(n110) );
  MUX21X1 U150 ( .IN1(n143), .IN2(n145), .S(SH[1]), .Q(n109) );
  MUX21X1 U151 ( .IN1(n142), .IN2(n144), .S(SH[1]), .Q(n108) );
  MUX21X1 U152 ( .IN1(n141), .IN2(n143), .S(SH[1]), .Q(n107) );
  MUX21X1 U153 ( .IN1(n140), .IN2(n142), .S(SH[1]), .Q(n106) );
  MUX21X1 U154 ( .IN1(n139), .IN2(n141), .S(SH[1]), .Q(n105) );
  MUX21X1 U155 ( .IN1(n138), .IN2(n140), .S(SH[1]), .Q(n104) );
  MUX21X1 U156 ( .IN1(n137), .IN2(n139), .S(SH[1]), .Q(n103) );
  MUX21X1 U157 ( .IN1(n136), .IN2(n138), .S(SH[1]), .Q(n102) );
  MUX21X1 U158 ( .IN1(n135), .IN2(n137), .S(SH[1]), .Q(n101) );
  MUX21X1 U159 ( .IN1(n134), .IN2(n136), .S(SH[1]), .Q(n100) );
  MUX21X1 U160 ( .IN1(n133), .IN2(n135), .S(SH[1]), .Q(n99) );
  MUX21X1 U161 ( .IN1(n132), .IN2(n134), .S(SH[1]), .Q(n98) );
  MUX21X1 U162 ( .IN1(n131), .IN2(n133), .S(SH[1]), .Q(n97) );
  MUX21X1 U165 ( .IN1(A[31]), .IN2(A[32]), .S(SH[0]), .Q(n162) );
  MUX21X1 U166 ( .IN1(A[30]), .IN2(A[31]), .S(SH[0]), .Q(n161) );
  MUX21X1 U167 ( .IN1(A[29]), .IN2(A[30]), .S(SH[0]), .Q(n160) );
  MUX21X1 U168 ( .IN1(A[28]), .IN2(A[29]), .S(SH[0]), .Q(n159) );
  MUX21X1 U169 ( .IN1(A[27]), .IN2(A[28]), .S(SH[0]), .Q(n158) );
  MUX21X1 U170 ( .IN1(A[26]), .IN2(A[27]), .S(SH[0]), .Q(n157) );
  MUX21X1 U171 ( .IN1(A[25]), .IN2(A[26]), .S(SH[0]), .Q(n156) );
  MUX21X1 U172 ( .IN1(A[24]), .IN2(A[25]), .S(SH[0]), .Q(n155) );
  MUX21X1 U173 ( .IN1(A[23]), .IN2(A[24]), .S(SH[0]), .Q(n154) );
  MUX21X1 U174 ( .IN1(A[22]), .IN2(A[23]), .S(SH[0]), .Q(n153) );
  MUX21X1 U175 ( .IN1(A[21]), .IN2(A[22]), .S(SH[0]), .Q(n152) );
  MUX21X1 U176 ( .IN1(A[20]), .IN2(A[21]), .S(SH[0]), .Q(n151) );
  MUX21X1 U177 ( .IN1(A[19]), .IN2(A[20]), .S(SH[0]), .Q(n150) );
  MUX21X1 U178 ( .IN1(A[18]), .IN2(A[19]), .S(SH[0]), .Q(n149) );
  MUX21X1 U179 ( .IN1(A[17]), .IN2(A[18]), .S(SH[0]), .Q(n148) );
  MUX21X1 U180 ( .IN1(A[16]), .IN2(A[17]), .S(SH[0]), .Q(n147) );
  MUX21X1 U181 ( .IN1(A[15]), .IN2(A[16]), .S(SH[0]), .Q(n146) );
  MUX21X1 U182 ( .IN1(A[14]), .IN2(A[15]), .S(SH[0]), .Q(n145) );
  MUX21X1 U183 ( .IN1(A[13]), .IN2(A[14]), .S(SH[0]), .Q(n144) );
  MUX21X1 U184 ( .IN1(A[12]), .IN2(A[13]), .S(SH[0]), .Q(n143) );
  MUX21X1 U185 ( .IN1(A[11]), .IN2(A[12]), .S(SH[0]), .Q(n142) );
  MUX21X1 U186 ( .IN1(A[10]), .IN2(A[11]), .S(SH[0]), .Q(n141) );
  MUX21X1 U187 ( .IN1(A[9]), .IN2(A[10]), .S(SH[0]), .Q(n140) );
  MUX21X1 U188 ( .IN1(A[8]), .IN2(A[9]), .S(SH[0]), .Q(n139) );
  MUX21X1 U189 ( .IN1(A[7]), .IN2(A[8]), .S(SH[0]), .Q(n138) );
  MUX21X1 U190 ( .IN1(A[6]), .IN2(A[7]), .S(SH[0]), .Q(n137) );
  MUX21X1 U191 ( .IN1(A[5]), .IN2(A[6]), .S(SH[0]), .Q(n136) );
  MUX21X1 U192 ( .IN1(A[4]), .IN2(A[5]), .S(SH[0]), .Q(n135) );
  MUX21X1 U193 ( .IN1(A[3]), .IN2(A[4]), .S(SH[0]), .Q(n134) );
  MUX21X1 U194 ( .IN1(A[2]), .IN2(A[3]), .S(SH[0]), .Q(n133) );
  MUX21X1 U195 ( .IN1(A[1]), .IN2(A[2]), .S(SH[0]), .Q(n132) );
  AND2X1 U196 ( .IN1(SH[0]), .IN2(A[1]), .Q(n131) );
  AND2X1 U200 ( .IN1(n56), .IN2(n1), .Q(B[31]) );
  AND2X1 U201 ( .IN1(n55), .IN2(n1), .Q(B[30]) );
  AND2X1 U202 ( .IN1(n54), .IN2(n1), .Q(B[29]) );
  AND2X1 U203 ( .IN1(n53), .IN2(n1), .Q(B[28]) );
  AND2X1 U204 ( .IN1(n52), .IN2(n1), .Q(B[27]) );
  AND2X1 U205 ( .IN1(n51), .IN2(n1), .Q(B[26]) );
  AND2X1 U206 ( .IN1(n50), .IN2(n1), .Q(B[25]) );
  AND2X1 U207 ( .IN1(n49), .IN2(n1), .Q(B[24]) );
  AND2X1 U208 ( .IN1(n48), .IN2(n1), .Q(B[23]) );
  AND2X1 U209 ( .IN1(n47), .IN2(n1), .Q(B[22]) );
  AND2X1 U210 ( .IN1(n46), .IN2(n1), .Q(B[21]) );
  AND2X1 U211 ( .IN1(n44), .IN2(n1), .Q(B[19]) );
  AND2X1 U212 ( .IN1(n43), .IN2(n1), .Q(B[18]) );
  AND2X1 U213 ( .IN1(n42), .IN2(n1), .Q(B[17]) );
  AND2X1 U214 ( .IN1(n45), .IN2(n1), .Q(B[20]) );
  AND2X1 U215 ( .IN1(n94), .IN2(n17), .Q(n57) );
  AND2X1 U216 ( .IN1(n93), .IN2(n17), .Q(n56) );
  AND2X1 U217 ( .IN1(n92), .IN2(n17), .Q(n55) );
  AND2X1 U218 ( .IN1(n91), .IN2(n17), .Q(n54) );
  AND2X1 U219 ( .IN1(n90), .IN2(n17), .Q(n53) );
  AND2X1 U220 ( .IN1(n89), .IN2(n17), .Q(n52) );
  AND2X1 U221 ( .IN1(n88), .IN2(n17), .Q(n51) );
  AND2X1 U222 ( .IN1(n87), .IN2(n17), .Q(n50) );
  AND2X1 U223 ( .IN1(n129), .IN2(n58), .Q(n94) );
  AND2X1 U224 ( .IN1(n128), .IN2(n58), .Q(n93) );
  AND2X1 U225 ( .IN1(n127), .IN2(n58), .Q(n92) );
  AND2X1 U226 ( .IN1(n126), .IN2(n58), .Q(n91) );
  AND2X1 U227 ( .IN1(n163), .IN2(n95), .Q(n129) );
  AND2X1 U228 ( .IN1(n162), .IN2(n95), .Q(n128) );
  AND2X1 U229 ( .IN1(n57), .IN2(n1), .Q(B[32]) );
  INVX0 U230 ( .INP(SH[4]), .ZN(n1) );
  INVX0 U231 ( .INP(SH[3]), .ZN(n17) );
  INVX0 U232 ( .INP(SH[2]), .ZN(n58) );
  INVX0 U233 ( .INP(SH[1]), .ZN(n95) );
  AND2X1 U234 ( .IN1(A[32]), .IN2(n130), .Q(n163) );
  INVX0 U235 ( .INP(SH[0]), .ZN(n130) );
endmodule


module thumb_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n2, n3, n5, n8, n9, n12, n13, n15, n17, n19, n21, n24, n28, n30, n32,
         n45, n46, n47, n48, n50, n51, n53, n55, n57, n59, n62, n64, n65, n67,
         n69, n74, n76, n78, n80, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604;

  XOR2X1 U83 ( .IN1(n98), .IN2(n97), .Q(product[31]) );
  XOR2X1 U84 ( .IN1(n128), .IN2(n158), .Q(n97) );
  FADDX1 U85 ( .A(n159), .B(n216), .CI(n99), .CO(n98), .S(product[30]) );
  FADDX1 U86 ( .A(n217), .B(n272), .CI(n100), .CO(n99), .S(product[29]) );
  FADDX1 U87 ( .A(n273), .B(n326), .CI(n101), .CO(n100), .S(product[28]) );
  FADDX1 U88 ( .A(n327), .B(n378), .CI(n102), .CO(n101), .S(product[27]) );
  FADDX1 U89 ( .A(n379), .B(n428), .CI(n103), .CO(n102), .S(product[26]) );
  FADDX1 U90 ( .A(n429), .B(n476), .CI(n104), .CO(n103), .S(product[25]) );
  FADDX1 U91 ( .A(n477), .B(n522), .CI(n105), .CO(n104), .S(product[24]) );
  FADDX1 U92 ( .A(n523), .B(n566), .CI(n106), .CO(n105), .S(product[23]) );
  FADDX1 U93 ( .A(n567), .B(n608), .CI(n107), .CO(n106), .S(product[22]) );
  FADDX1 U94 ( .A(n609), .B(n648), .CI(n108), .CO(n107), .S(product[21]) );
  FADDX1 U95 ( .A(n649), .B(n686), .CI(n109), .CO(n108), .S(product[20]) );
  FADDX1 U96 ( .A(n687), .B(n722), .CI(n110), .CO(n109), .S(product[19]) );
  FADDX1 U97 ( .A(n723), .B(n756), .CI(n111), .CO(n110), .S(product[18]) );
  FADDX1 U98 ( .A(n757), .B(n788), .CI(n112), .CO(n111), .S(product[17]) );
  FADDX1 U99 ( .A(n789), .B(n818), .CI(n113), .CO(n112), .S(product[16]) );
  FADDX1 U100 ( .A(n819), .B(n846), .CI(n114), .CO(n113), .S(product[15]) );
  FADDX1 U101 ( .A(n847), .B(n872), .CI(n115), .CO(n114), .S(product[14]) );
  FADDX1 U102 ( .A(n873), .B(n896), .CI(n116), .CO(n115), .S(product[13]) );
  FADDX1 U103 ( .A(n897), .B(n918), .CI(n117), .CO(n116), .S(product[12]) );
  FADDX1 U104 ( .A(n919), .B(n938), .CI(n118), .CO(n117), .S(product[11]) );
  FADDX1 U105 ( .A(n939), .B(n956), .CI(n119), .CO(n118), .S(product[10]) );
  FADDX1 U106 ( .A(n957), .B(n972), .CI(n120), .CO(n119), .S(product[9]) );
  FADDX1 U107 ( .A(n973), .B(n986), .CI(n121), .CO(n120), .S(product[8]) );
  FADDX1 U108 ( .A(n987), .B(n998), .CI(n122), .CO(n121), .S(product[7]) );
  FADDX1 U109 ( .A(n999), .B(n1008), .CI(n123), .CO(n122), .S(product[6]) );
  FADDX1 U110 ( .A(n1009), .B(n1016), .CI(n124), .CO(n123), .S(product[5]) );
  FADDX1 U111 ( .A(n1017), .B(n1022), .CI(n125), .CO(n124), .S(product[4]) );
  FADDX1 U112 ( .A(n1023), .B(n1026), .CI(n126), .CO(n125), .S(product[3]) );
  FADDX1 U113 ( .A(n1027), .B(n1492), .CI(n127), .CO(n126), .S(product[2]) );
  HADDX1 U114 ( .A0(n1523), .B0(n1554), .C1(n127), .SO(product[1]) );
  XOR3X1 U115 ( .IN1(n130), .IN2(n160), .IN3(n129), .Q(n128) );
  XOR3X1 U116 ( .IN1(n132), .IN2(n162), .IN3(n131), .Q(n129) );
  XOR3X1 U117 ( .IN1(n164), .IN2(n134), .IN3(n133), .Q(n130) );
  XOR3X1 U118 ( .IN1(n136), .IN2(n166), .IN3(n135), .Q(n131) );
  XOR3X1 U119 ( .IN1(n137), .IN2(n170), .IN3(n168), .Q(n132) );
  XOR3X1 U120 ( .IN1(n139), .IN2(n141), .IN3(n138), .Q(n133) );
  XOR3X1 U121 ( .IN1(n140), .IN2(n172), .IN3(n142), .Q(n134) );
  XOR3X1 U122 ( .IN1(n176), .IN2(n178), .IN3(n174), .Q(n135) );
  XOR3X1 U123 ( .IN1(n144), .IN2(n143), .IN3(n180), .Q(n136) );
  XOR3X1 U124 ( .IN1(n146), .IN2(n184), .IN3(n145), .Q(n137) );
  XOR3X1 U125 ( .IN1(n188), .IN2(n186), .IN3(n182), .Q(n138) );
  XOR3X1 U126 ( .IN1(n192), .IN2(n148), .IN3(n190), .Q(n139) );
  XOR3X1 U127 ( .IN1(n150), .IN2(n153), .IN3(n154), .Q(n140) );
  XOR3X1 U128 ( .IN1(n151), .IN2(n152), .IN3(n149), .Q(n141) );
  XOR3X1 U129 ( .IN1(n156), .IN2(n147), .IN3(n155), .Q(n142) );
  XOR3X1 U130 ( .IN1(n202), .IN2(n206), .IN3(n194), .Q(n143) );
  XOR3X1 U131 ( .IN1(n200), .IN2(n204), .IN3(n208), .Q(n144) );
  XOR3X1 U132 ( .IN1(n210), .IN2(n196), .IN3(n198), .Q(n145) );
  XOR3X1 U133 ( .IN1(n214), .IN2(n157), .IN3(n212), .Q(n146) );
  XOR3X1 U134 ( .IN1(n1218), .IN2(n1259), .IN3(n1238), .Q(n147) );
  XOR3X1 U135 ( .IN1(n1106), .IN2(n1281), .IN3(n1199), .Q(n148) );
  XOR3X1 U136 ( .IN1(n1073), .IN2(n1304), .IN3(n1094), .Q(n149) );
  XOR3X1 U137 ( .IN1(n1056), .IN2(n1328), .IN3(n1064), .Q(n150) );
  XOR3X1 U138 ( .IN1(n1379), .IN2(n1083), .IN3(n1353), .Q(n151) );
  XOR3X1 U139 ( .IN1(n1406), .IN2(n1119), .IN3(n1049), .Q(n152) );
  XOR3X1 U140 ( .IN1(n1043), .IN2(n1164), .IN3(n1434), .Q(n153) );
  XOR3X1 U141 ( .IN1(n1463), .IN2(n1133), .IN3(n1038), .Q(n154) );
  XOR3X1 U142 ( .IN1(n1493), .IN2(n1148), .IN3(n1034), .Q(n155) );
  XOR3X1 U143 ( .IN1(n1524), .IN2(n1181), .IN3(n1031), .Q(n156) );
  XOR2X1 U144 ( .IN1(n1028), .IN2(n1029), .Q(n157) );
  FADDX1 U145 ( .A(n218), .B(n163), .CI(n161), .CO(n158), .S(n159) );
  FADDX1 U146 ( .A(n165), .B(n222), .CI(n220), .CO(n160), .S(n161) );
  FADDX1 U147 ( .A(n169), .B(n167), .CI(n224), .CO(n162), .S(n163) );
  FADDX1 U148 ( .A(n171), .B(n228), .CI(n226), .CO(n164), .S(n165) );
  FADDX1 U149 ( .A(n179), .B(n230), .CI(n175), .CO(n166), .S(n167) );
  FADDX1 U150 ( .A(n177), .B(n232), .CI(n173), .CO(n168), .S(n169) );
  FADDX1 U151 ( .A(n236), .B(n181), .CI(n234), .CO(n170), .S(n171) );
  FADDX1 U152 ( .A(n191), .B(n238), .CI(n185), .CO(n172), .S(n173) );
  FADDX1 U153 ( .A(n240), .B(n193), .CI(n183), .CO(n174), .S(n175) );
  FADDX1 U154 ( .A(n244), .B(n246), .CI(n189), .CO(n176), .S(n177) );
  FADDX1 U155 ( .A(n242), .B(n248), .CI(n187), .CO(n178), .S(n179) );
  FADDX1 U156 ( .A(n195), .B(n199), .CI(n250), .CO(n180), .S(n181) );
  FADDX1 U157 ( .A(n201), .B(n203), .CI(n213), .CO(n182), .S(n183) );
  FADDX1 U158 ( .A(n209), .B(n266), .CI(n205), .CO(n184), .S(n185) );
  FADDX1 U159 ( .A(n264), .B(n260), .CI(n207), .CO(n186), .S(n187) );
  FADDX1 U160 ( .A(n258), .B(n262), .CI(n211), .CO(n188), .S(n189) );
  FADDX1 U161 ( .A(n268), .B(n252), .CI(n197), .CO(n190), .S(n191) );
  FADDX1 U162 ( .A(n254), .B(n270), .CI(n256), .CO(n192), .S(n193) );
  FADDX1 U163 ( .A(n1260), .B(n1282), .CI(n215), .CO(n194), .S(n195) );
  FADDX1 U164 ( .A(n1219), .B(n1305), .CI(n1239), .CO(n196), .S(n197) );
  FADDX1 U165 ( .A(n1120), .B(n1329), .CI(n1182), .CO(n198), .S(n199) );
  FADDX1 U166 ( .A(n1084), .B(n1354), .CI(n1095), .CO(n200), .S(n201) );
  FADDX1 U167 ( .A(n1065), .B(n1057), .CI(n1074), .CO(n202), .S(n203) );
  FADDX1 U168 ( .A(n1050), .B(n1107), .CI(n1380), .CO(n204), .S(n205) );
  FADDX1 U169 ( .A(n1435), .B(n1165), .CI(n1407), .CO(n206), .S(n207) );
  FADDX1 U170 ( .A(n1464), .B(n1134), .CI(n1044), .CO(n208), .S(n209) );
  FADDX1 U171 ( .A(n1039), .B(n1149), .CI(n1494), .CO(n210), .S(n211) );
  FADDX1 U172 ( .A(n1035), .B(n1200), .CI(n1525), .CO(n212), .S(n213) );
  HADDX1 U173 ( .A0(n1032), .B0(n1030), .C1(n214), .SO(n215) );
  FADDX1 U174 ( .A(n274), .B(n221), .CI(n219), .CO(n216), .S(n217) );
  FADDX1 U175 ( .A(n223), .B(n278), .CI(n276), .CO(n218), .S(n219) );
  FADDX1 U176 ( .A(n227), .B(n280), .CI(n225), .CO(n220), .S(n221) );
  FADDX1 U177 ( .A(n229), .B(n284), .CI(n282), .CO(n222), .S(n223) );
  FADDX1 U178 ( .A(n231), .B(n286), .CI(n233), .CO(n224), .S(n225) );
  FADDX1 U179 ( .A(n288), .B(n290), .CI(n235), .CO(n226), .S(n227) );
  FADDX1 U180 ( .A(n292), .B(n294), .CI(n237), .CO(n228), .S(n229) );
  FADDX1 U181 ( .A(n243), .B(n296), .CI(n241), .CO(n230), .S(n231) );
  FADDX1 U182 ( .A(n245), .B(n247), .CI(n239), .CO(n232), .S(n233) );
  FADDX1 U183 ( .A(n300), .B(n302), .CI(n249), .CO(n234), .S(n235) );
  FADDX1 U184 ( .A(n304), .B(n251), .CI(n298), .CO(n236), .S(n237) );
  FADDX1 U185 ( .A(n257), .B(n259), .CI(n269), .CO(n238), .S(n239) );
  FADDX1 U186 ( .A(n263), .B(n312), .CI(n261), .CO(n240), .S(n241) );
  FADDX1 U187 ( .A(n316), .B(n314), .CI(n265), .CO(n242), .S(n243) );
  FADDX1 U188 ( .A(n318), .B(n306), .CI(n267), .CO(n244), .S(n245) );
  FADDX1 U189 ( .A(n320), .B(n310), .CI(n255), .CO(n246), .S(n247) );
  FADDX1 U190 ( .A(n322), .B(n308), .CI(n253), .CO(n248), .S(n249) );
  FADDX1 U191 ( .A(n271), .B(n1306), .CI(n324), .CO(n250), .S(n251) );
  FADDX1 U192 ( .A(n1330), .B(n1355), .CI(n1283), .CO(n252), .S(n253) );
  FADDX1 U193 ( .A(n1183), .B(n1381), .CI(n1261), .CO(n254), .S(n255) );
  FADDX1 U194 ( .A(n1121), .B(n1408), .CI(n1135), .CO(n256), .S(n257) );
  FADDX1 U195 ( .A(n1096), .B(n1436), .CI(n1108), .CO(n258), .S(n259) );
  FADDX1 U196 ( .A(n1085), .B(n1240), .CI(n1465), .CO(n260), .S(n261) );
  FADDX1 U197 ( .A(n1066), .B(n1220), .CI(n1075), .CO(n262), .S(n263) );
  FADDX1 U198 ( .A(n1051), .B(n1166), .CI(n1058), .CO(n264), .S(n265) );
  FADDX1 U199 ( .A(n1040), .B(n1150), .CI(n1045), .CO(n266), .S(n267) );
  FADDX1 U200 ( .A(n1526), .B(n1201), .CI(n1495), .CO(n268), .S(n269) );
  HADDX1 U201 ( .A0(n1036), .B0(n1033), .C1(n270), .SO(n271) );
  FADDX1 U202 ( .A(n328), .B(n277), .CI(n275), .CO(n272), .S(n273) );
  FADDX1 U203 ( .A(n279), .B(n332), .CI(n330), .CO(n274), .S(n275) );
  FADDX1 U204 ( .A(n283), .B(n334), .CI(n281), .CO(n276), .S(n277) );
  FADDX1 U205 ( .A(n285), .B(n338), .CI(n336), .CO(n278), .S(n279) );
  FADDX1 U206 ( .A(n289), .B(n340), .CI(n287), .CO(n280), .S(n281) );
  FADDX1 U207 ( .A(n342), .B(n344), .CI(n291), .CO(n282), .S(n283) );
  FADDX1 U208 ( .A(n346), .B(n297), .CI(n293), .CO(n284), .S(n285) );
  FADDX1 U209 ( .A(n301), .B(n348), .CI(n295), .CO(n286), .S(n287) );
  FADDX1 U210 ( .A(n352), .B(n354), .CI(n299), .CO(n288), .S(n289) );
  FADDX1 U211 ( .A(n350), .B(n356), .CI(n303), .CO(n290), .S(n291) );
  FADDX1 U212 ( .A(n358), .B(n313), .CI(n305), .CO(n292), .S(n293) );
  FADDX1 U213 ( .A(n309), .B(n321), .CI(n311), .CO(n294), .S(n295) );
  FADDX1 U214 ( .A(n319), .B(n368), .CI(n315), .CO(n296), .S(n297) );
  FADDX1 U215 ( .A(n362), .B(n364), .CI(n317), .CO(n298), .S(n299) );
  FADDX1 U216 ( .A(n370), .B(n366), .CI(n323), .CO(n300), .S(n301) );
  FADDX1 U217 ( .A(n372), .B(n360), .CI(n307), .CO(n302), .S(n303) );
  FADDX1 U218 ( .A(n376), .B(n325), .CI(n374), .CO(n304), .S(n305) );
  FADDX1 U219 ( .A(n1307), .B(n1331), .CI(n1284), .CO(n306), .S(n307) );
  FADDX1 U220 ( .A(n1151), .B(n1356), .CI(n1262), .CO(n308), .S(n309) );
  FADDX1 U221 ( .A(n1122), .B(n1382), .CI(n1136), .CO(n310), .S(n311) );
  FADDX1 U222 ( .A(n1097), .B(n1409), .CI(n1109), .CO(n312), .S(n313) );
  FADDX1 U223 ( .A(n1466), .B(n1241), .CI(n1437), .CO(n314), .S(n315) );
  FADDX1 U224 ( .A(n1076), .B(n1167), .CI(n1086), .CO(n316), .S(n317) );
  FADDX1 U225 ( .A(n1067), .B(n1202), .CI(n1496), .CO(n318), .S(n319) );
  FADDX1 U226 ( .A(n1059), .B(n1184), .CI(n1527), .CO(n320), .S(n321) );
  FADDX1 U227 ( .A(n1046), .B(n1221), .CI(n1052), .CO(n322), .S(n323) );
  HADDX1 U228 ( .A0(n1041), .B0(n1037), .C1(n324), .SO(n325) );
  FADDX1 U229 ( .A(n380), .B(n331), .CI(n329), .CO(n326), .S(n327) );
  FADDX1 U230 ( .A(n333), .B(n384), .CI(n382), .CO(n328), .S(n329) );
  FADDX1 U231 ( .A(n386), .B(n337), .CI(n335), .CO(n330), .S(n331) );
  FADDX1 U232 ( .A(n339), .B(n390), .CI(n388), .CO(n332), .S(n333) );
  FADDX1 U233 ( .A(n343), .B(n392), .CI(n341), .CO(n334), .S(n335) );
  FADDX1 U234 ( .A(n394), .B(n396), .CI(n345), .CO(n336), .S(n337) );
  FADDX1 U235 ( .A(n355), .B(n351), .CI(n347), .CO(n338), .S(n339) );
  FADDX1 U236 ( .A(n398), .B(n357), .CI(n349), .CO(n340), .S(n341) );
  FADDX1 U237 ( .A(n404), .B(n406), .CI(n353), .CO(n342), .S(n343) );
  FADDX1 U238 ( .A(n402), .B(n408), .CI(n400), .CO(n344), .S(n345) );
  FADDX1 U239 ( .A(n369), .B(n363), .CI(n359), .CO(n346), .S(n347) );
  FADDX1 U240 ( .A(n365), .B(n373), .CI(n367), .CO(n348), .S(n349) );
  FADDX1 U241 ( .A(n418), .B(n416), .CI(n375), .CO(n350), .S(n351) );
  FADDX1 U242 ( .A(n422), .B(n420), .CI(n371), .CO(n352), .S(n353) );
  FADDX1 U243 ( .A(n424), .B(n410), .CI(n361), .CO(n354), .S(n355) );
  FADDX1 U244 ( .A(n412), .B(n426), .CI(n414), .CO(n356), .S(n357) );
  FADDX1 U245 ( .A(n1263), .B(n1242), .CI(n377), .CO(n358), .S(n359) );
  FADDX1 U246 ( .A(n1168), .B(n1285), .CI(n1203), .CO(n360), .S(n361) );
  FADDX1 U247 ( .A(n1098), .B(n1308), .CI(n1110), .CO(n362), .S(n363) );
  FADDX1 U248 ( .A(n1077), .B(n1332), .CI(n1087), .CO(n364), .S(n365) );
  FADDX1 U249 ( .A(n1068), .B(n1137), .CI(n1357), .CO(n366), .S(n367) );
  FADDX1 U250 ( .A(n1383), .B(n1123), .CI(n1060), .CO(n368), .S(n369) );
  FADDX1 U251 ( .A(n1438), .B(n1152), .CI(n1410), .CO(n370), .S(n371) );
  FADDX1 U252 ( .A(n1497), .B(n1185), .CI(n1467), .CO(n372), .S(n373) );
  FADDX1 U253 ( .A(n1528), .B(n1222), .CI(n1053), .CO(n374), .S(n375) );
  HADDX1 U254 ( .A0(n1047), .B0(n1042), .C1(n376), .SO(n377) );
  FADDX1 U255 ( .A(n430), .B(n383), .CI(n381), .CO(n378), .S(n379) );
  FADDX1 U256 ( .A(n385), .B(n434), .CI(n432), .CO(n380), .S(n381) );
  FADDX1 U257 ( .A(n436), .B(n389), .CI(n387), .CO(n382), .S(n383) );
  FADDX1 U258 ( .A(n393), .B(n440), .CI(n438), .CO(n384), .S(n385) );
  FADDX1 U259 ( .A(n395), .B(n442), .CI(n391), .CO(n386), .S(n387) );
  FADDX1 U260 ( .A(n397), .B(n446), .CI(n444), .CO(n388), .S(n389) );
  FADDX1 U261 ( .A(n403), .B(n448), .CI(n399), .CO(n390), .S(n391) );
  FADDX1 U262 ( .A(n407), .B(n454), .CI(n401), .CO(n392), .S(n393) );
  FADDX1 U263 ( .A(n452), .B(n450), .CI(n405), .CO(n394), .S(n395) );
  FADDX1 U264 ( .A(n409), .B(n419), .CI(n456), .CO(n396), .S(n397) );
  FADDX1 U265 ( .A(n415), .B(n423), .CI(n417), .CO(n398), .S(n399) );
  FADDX1 U266 ( .A(n468), .B(n466), .CI(n421), .CO(n400), .S(n401) );
  FADDX1 U267 ( .A(n470), .B(n464), .CI(n425), .CO(n402), .S(n403) );
  FADDX1 U268 ( .A(n472), .B(n462), .CI(n413), .CO(n404), .S(n405) );
  FADDX1 U269 ( .A(n458), .B(n460), .CI(n411), .CO(n406), .S(n407) );
  FADDX1 U270 ( .A(n427), .B(n1358), .CI(n474), .CO(n408), .S(n409) );
  FADDX1 U271 ( .A(n1309), .B(n1384), .CI(n1333), .CO(n410), .S(n411) );
  FADDX1 U272 ( .A(n1169), .B(n1411), .CI(n1286), .CO(n412), .S(n413) );
  FADDX1 U273 ( .A(n1138), .B(n1439), .CI(n1153), .CO(n414), .S(n415) );
  FADDX1 U274 ( .A(n1124), .B(n1264), .CI(n1468), .CO(n416), .S(n417) );
  FADDX1 U275 ( .A(n1099), .B(n1223), .CI(n1111), .CO(n418), .S(n419) );
  FADDX1 U276 ( .A(n1078), .B(n1204), .CI(n1088), .CO(n420), .S(n421) );
  FADDX1 U277 ( .A(n1498), .B(n1186), .CI(n1069), .CO(n422), .S(n423) );
  FADDX1 U278 ( .A(n1061), .B(n1243), .CI(n1529), .CO(n424), .S(n425) );
  HADDX1 U279 ( .A0(n1054), .B0(n1048), .C1(n426), .SO(n427) );
  FADDX1 U280 ( .A(n478), .B(n433), .CI(n431), .CO(n428), .S(n429) );
  FADDX1 U281 ( .A(n435), .B(n437), .CI(n480), .CO(n430), .S(n431) );
  FADDX1 U282 ( .A(n484), .B(n439), .CI(n482), .CO(n432), .S(n433) );
  FADDX1 U283 ( .A(n441), .B(n443), .CI(n486), .CO(n434), .S(n435) );
  FADDX1 U284 ( .A(n445), .B(n490), .CI(n488), .CO(n436), .S(n437) );
  FADDX1 U285 ( .A(n447), .B(n494), .CI(n492), .CO(n438), .S(n439) );
  FADDX1 U286 ( .A(n451), .B(n496), .CI(n449), .CO(n440), .S(n441) );
  FADDX1 U287 ( .A(n455), .B(n498), .CI(n453), .CO(n442), .S(n443) );
  FADDX1 U288 ( .A(n500), .B(n457), .CI(n502), .CO(n444), .S(n445) );
  FADDX1 U289 ( .A(n467), .B(n461), .CI(n504), .CO(n446), .S(n447) );
  FADDX1 U290 ( .A(n463), .B(n471), .CI(n465), .CO(n448), .S(n449) );
  FADDX1 U291 ( .A(n510), .B(n508), .CI(n473), .CO(n450), .S(n451) );
  FADDX1 U292 ( .A(n514), .B(n512), .CI(n469), .CO(n452), .S(n453) );
  FADDX1 U293 ( .A(n516), .B(n506), .CI(n459), .CO(n454), .S(n455) );
  FADDX1 U294 ( .A(n520), .B(n475), .CI(n518), .CO(n456), .S(n457) );
  FADDX1 U295 ( .A(n1265), .B(n1310), .CI(n1287), .CO(n458), .S(n459) );
  FADDX1 U296 ( .A(n1205), .B(n1334), .CI(n1224), .CO(n460), .S(n461) );
  FADDX1 U297 ( .A(n1125), .B(n1359), .CI(n1170), .CO(n462), .S(n463) );
  FADDX1 U298 ( .A(n1100), .B(n1089), .CI(n1112), .CO(n464), .S(n465) );
  FADDX1 U299 ( .A(n1070), .B(n1139), .CI(n1079), .CO(n466), .S(n467) );
  FADDX1 U300 ( .A(n1412), .B(n1154), .CI(n1385), .CO(n468), .S(n469) );
  FADDX1 U301 ( .A(n1469), .B(n1187), .CI(n1440), .CO(n470), .S(n471) );
  FADDX1 U302 ( .A(n1530), .B(n1244), .CI(n1499), .CO(n472), .S(n473) );
  HADDX1 U303 ( .A0(n1062), .B0(n1055), .C1(n474), .SO(n475) );
  FADDX1 U304 ( .A(n524), .B(n481), .CI(n479), .CO(n476), .S(n477) );
  FADDX1 U305 ( .A(n483), .B(n528), .CI(n526), .CO(n478), .S(n479) );
  FADDX1 U306 ( .A(n530), .B(n487), .CI(n485), .CO(n480), .S(n481) );
  FADDX1 U307 ( .A(n491), .B(n534), .CI(n489), .CO(n482), .S(n483) );
  FADDX1 U308 ( .A(n536), .B(n493), .CI(n532), .CO(n484), .S(n485) );
  FADDX1 U309 ( .A(n497), .B(n501), .CI(n538), .CO(n486), .S(n487) );
  FADDX1 U310 ( .A(n540), .B(n503), .CI(n495), .CO(n488), .S(n489) );
  FADDX1 U311 ( .A(n542), .B(n544), .CI(n499), .CO(n490), .S(n491) );
  FADDX1 U312 ( .A(n548), .B(n505), .CI(n546), .CO(n492), .S(n493) );
  FADDX1 U313 ( .A(n509), .B(n519), .CI(n507), .CO(n494), .S(n495) );
  FADDX1 U314 ( .A(n513), .B(n556), .CI(n511), .CO(n496), .S(n497) );
  FADDX1 U315 ( .A(n560), .B(n558), .CI(n515), .CO(n498), .S(n499) );
  FADDX1 U316 ( .A(n562), .B(n554), .CI(n517), .CO(n500), .S(n501) );
  FADDX1 U317 ( .A(n552), .B(n564), .CI(n550), .CO(n502), .S(n503) );
  FADDX1 U318 ( .A(n1245), .B(n1288), .CI(n521), .CO(n504), .S(n505) );
  FADDX1 U319 ( .A(n1188), .B(n1311), .CI(n1225), .CO(n506), .S(n507) );
  FADDX1 U320 ( .A(n1126), .B(n1335), .CI(n1140), .CO(n508), .S(n509) );
  FADDX1 U321 ( .A(n1101), .B(n1360), .CI(n1113), .CO(n510), .S(n511) );
  FADDX1 U322 ( .A(n1386), .B(n1155), .CI(n1090), .CO(n512), .S(n513) );
  FADDX1 U323 ( .A(n1441), .B(n1171), .CI(n1413), .CO(n514), .S(n515) );
  FADDX1 U324 ( .A(n1080), .B(n1206), .CI(n1470), .CO(n516), .S(n517) );
  FADDX1 U325 ( .A(n1531), .B(n1266), .CI(n1500), .CO(n518), .S(n519) );
  HADDX1 U326 ( .A0(n1071), .B0(n1063), .C1(n520), .SO(n521) );
  FADDX1 U327 ( .A(n568), .B(n527), .CI(n525), .CO(n522), .S(n523) );
  FADDX1 U328 ( .A(n529), .B(n572), .CI(n570), .CO(n524), .S(n525) );
  FADDX1 U329 ( .A(n574), .B(n533), .CI(n531), .CO(n526), .S(n527) );
  FADDX1 U330 ( .A(n576), .B(n537), .CI(n535), .CO(n528), .S(n529) );
  FADDX1 U331 ( .A(n580), .B(n539), .CI(n578), .CO(n530), .S(n531) );
  FADDX1 U332 ( .A(n545), .B(n584), .CI(n582), .CO(n532), .S(n533) );
  FADDX1 U333 ( .A(n543), .B(n547), .CI(n541), .CO(n534), .S(n535) );
  FADDX1 U334 ( .A(n586), .B(n590), .CI(n588), .CO(n536), .S(n537) );
  FADDX1 U335 ( .A(n555), .B(n559), .CI(n549), .CO(n538), .S(n539) );
  FADDX1 U336 ( .A(n561), .B(n596), .CI(n553), .CO(n540), .S(n541) );
  FADDX1 U337 ( .A(n600), .B(n598), .CI(n557), .CO(n542), .S(n543) );
  FADDX1 U338 ( .A(n602), .B(n592), .CI(n563), .CO(n544), .S(n545) );
  FADDX1 U339 ( .A(n604), .B(n594), .CI(n551), .CO(n546), .S(n547) );
  FADDX1 U340 ( .A(n565), .B(n1312), .CI(n606), .CO(n548), .S(n549) );
  FADDX1 U341 ( .A(n1361), .B(n1387), .CI(n1336), .CO(n550), .S(n551) );
  FADDX1 U342 ( .A(n1189), .B(n1414), .CI(n1289), .CO(n552), .S(n553) );
  FADDX1 U343 ( .A(n1156), .B(n1442), .CI(n1172), .CO(n554), .S(n555) );
  FADDX1 U344 ( .A(n1127), .B(n1246), .CI(n1141), .CO(n556), .S(n557) );
  FADDX1 U345 ( .A(n1471), .B(n1207), .CI(n1114), .CO(n558), .S(n559) );
  FADDX1 U346 ( .A(n1501), .B(n1226), .CI(n1102), .CO(n560), .S(n561) );
  FADDX1 U347 ( .A(n1532), .B(n1267), .CI(n1091), .CO(n562), .S(n563) );
  HADDX1 U348 ( .A0(n1081), .B0(n1072), .C1(n564), .SO(n565) );
  FADDX1 U349 ( .A(n610), .B(n571), .CI(n569), .CO(n566), .S(n567) );
  FADDX1 U350 ( .A(n573), .B(n614), .CI(n612), .CO(n568), .S(n569) );
  FADDX1 U351 ( .A(n616), .B(n577), .CI(n575), .CO(n570), .S(n571) );
  FADDX1 U352 ( .A(n618), .B(n581), .CI(n579), .CO(n572), .S(n573) );
  FADDX1 U353 ( .A(n622), .B(n585), .CI(n620), .CO(n574), .S(n575) );
  FADDX1 U354 ( .A(n589), .B(n624), .CI(n583), .CO(n576), .S(n577) );
  FADDX1 U355 ( .A(n626), .B(n628), .CI(n587), .CO(n578), .S(n579) );
  FADDX1 U356 ( .A(n591), .B(n632), .CI(n630), .CO(n580), .S(n581) );
  FADDX1 U357 ( .A(n593), .B(n597), .CI(n599), .CO(n582), .S(n583) );
  FADDX1 U358 ( .A(n595), .B(n636), .CI(n603), .CO(n584), .S(n585) );
  FADDX1 U359 ( .A(n640), .B(n638), .CI(n601), .CO(n586), .S(n587) );
  FADDX1 U360 ( .A(n642), .B(n634), .CI(n605), .CO(n588), .S(n589) );
  FADDX1 U361 ( .A(n646), .B(n607), .CI(n644), .CO(n590), .S(n591) );
  FADDX1 U362 ( .A(n1313), .B(n1290), .CI(n1337), .CO(n592), .S(n593) );
  FADDX1 U363 ( .A(n1173), .B(n1362), .CI(n1208), .CO(n594), .S(n595) );
  FADDX1 U364 ( .A(n1142), .B(n1388), .CI(n1157), .CO(n596), .S(n597) );
  FADDX1 U365 ( .A(n1128), .B(n1190), .CI(n1415), .CO(n598), .S(n599) );
  FADDX1 U366 ( .A(n1472), .B(n1247), .CI(n1443), .CO(n600), .S(n601) );
  FADDX1 U367 ( .A(n1115), .B(n1227), .CI(n1502), .CO(n602), .S(n603) );
  FADDX1 U368 ( .A(n1533), .B(n1268), .CI(n1103), .CO(n604), .S(n605) );
  HADDX1 U369 ( .A0(n1092), .B0(n1082), .C1(n606), .SO(n607) );
  FADDX1 U370 ( .A(n650), .B(n613), .CI(n611), .CO(n608), .S(n609) );
  FADDX1 U371 ( .A(n652), .B(n654), .CI(n615), .CO(n610), .S(n611) );
  FADDX1 U372 ( .A(n619), .B(n621), .CI(n617), .CO(n612), .S(n613) );
  FADDX1 U373 ( .A(n658), .B(n660), .CI(n656), .CO(n614), .S(n615) );
  FADDX1 U374 ( .A(n625), .B(n662), .CI(n623), .CO(n616), .S(n617) );
  FADDX1 U375 ( .A(n631), .B(n666), .CI(n629), .CO(n618), .S(n619) );
  FADDX1 U376 ( .A(n664), .B(n668), .CI(n627), .CO(n620), .S(n621) );
  FADDX1 U377 ( .A(n633), .B(n641), .CI(n670), .CO(n622), .S(n623) );
  FADDX1 U378 ( .A(n635), .B(n645), .CI(n637), .CO(n624), .S(n625) );
  FADDX1 U379 ( .A(n682), .B(n680), .CI(n639), .CO(n626), .S(n627) );
  FADDX1 U380 ( .A(n678), .B(n676), .CI(n643), .CO(n628), .S(n629) );
  FADDX1 U381 ( .A(n674), .B(n684), .CI(n672), .CO(n630), .S(n631) );
  FADDX1 U382 ( .A(n1314), .B(n1338), .CI(n647), .CO(n632), .S(n633) );
  FADDX1 U383 ( .A(n1191), .B(n1363), .CI(n1209), .CO(n634), .S(n635) );
  FADDX1 U384 ( .A(n1158), .B(n1389), .CI(n1174), .CO(n636), .S(n637) );
  FADDX1 U385 ( .A(n1444), .B(n1269), .CI(n1416), .CO(n638), .S(n639) );
  FADDX1 U386 ( .A(n1473), .B(n1228), .CI(n1143), .CO(n640), .S(n641) );
  FADDX1 U387 ( .A(n1129), .B(n1248), .CI(n1503), .CO(n642), .S(n643) );
  FADDX1 U388 ( .A(n1534), .B(n1291), .CI(n1116), .CO(n644), .S(n645) );
  HADDX1 U389 ( .A0(n1104), .B0(n1093), .C1(n646), .SO(n647) );
  FADDX1 U390 ( .A(n688), .B(n653), .CI(n651), .CO(n648), .S(n649) );
  FADDX1 U391 ( .A(n655), .B(n692), .CI(n690), .CO(n650), .S(n651) );
  FADDX1 U392 ( .A(n659), .B(n694), .CI(n657), .CO(n652), .S(n653) );
  FADDX1 U393 ( .A(n661), .B(n698), .CI(n696), .CO(n654), .S(n655) );
  FADDX1 U394 ( .A(n667), .B(n700), .CI(n663), .CO(n656), .S(n657) );
  FADDX1 U395 ( .A(n665), .B(n702), .CI(n669), .CO(n658), .S(n659) );
  FADDX1 U396 ( .A(n706), .B(n671), .CI(n704), .CO(n660), .S(n661) );
  FADDX1 U397 ( .A(n675), .B(n677), .CI(n679), .CO(n662), .S(n663) );
  FADDX1 U398 ( .A(n714), .B(n712), .CI(n681), .CO(n664), .S(n665) );
  FADDX1 U399 ( .A(n716), .B(n708), .CI(n683), .CO(n666), .S(n667) );
  FADDX1 U400 ( .A(n718), .B(n710), .CI(n673), .CO(n668), .S(n669) );
  FADDX1 U401 ( .A(n685), .B(n1390), .CI(n720), .CO(n670), .S(n671) );
  FADDX1 U402 ( .A(n1339), .B(n1417), .CI(n1364), .CO(n672), .S(n673) );
  FADDX1 U403 ( .A(n1210), .B(n1445), .CI(n1315), .CO(n674), .S(n675) );
  FADDX1 U404 ( .A(n1175), .B(n1249), .CI(n1192), .CO(n676), .S(n677) );
  FADDX1 U405 ( .A(n1159), .B(n1270), .CI(n1474), .CO(n678), .S(n679) );
  FADDX1 U406 ( .A(n1130), .B(n1229), .CI(n1144), .CO(n680), .S(n681) );
  FADDX1 U407 ( .A(n1535), .B(n1292), .CI(n1504), .CO(n682), .S(n683) );
  HADDX1 U408 ( .A0(n1117), .B0(n1105), .C1(n684), .SO(n685) );
  FADDX1 U409 ( .A(n724), .B(n691), .CI(n689), .CO(n686), .S(n687) );
  FADDX1 U410 ( .A(n693), .B(n728), .CI(n726), .CO(n688), .S(n689) );
  FADDX1 U411 ( .A(n697), .B(n730), .CI(n695), .CO(n690), .S(n691) );
  FADDX1 U412 ( .A(n699), .B(n734), .CI(n732), .CO(n692), .S(n693) );
  FADDX1 U413 ( .A(n703), .B(n736), .CI(n701), .CO(n694), .S(n695) );
  FADDX1 U414 ( .A(n738), .B(n740), .CI(n705), .CO(n696), .S(n697) );
  FADDX1 U415 ( .A(n742), .B(n709), .CI(n707), .CO(n698), .S(n699) );
  FADDX1 U416 ( .A(n711), .B(n715), .CI(n717), .CO(n700), .S(n701) );
  FADDX1 U417 ( .A(n748), .B(n746), .CI(n713), .CO(n702), .S(n703) );
  FADDX1 U418 ( .A(n750), .B(n744), .CI(n719), .CO(n704), .S(n705) );
  FADDX1 U419 ( .A(n754), .B(n721), .CI(n752), .CO(n706), .S(n707) );
  FADDX1 U420 ( .A(n1293), .B(n1391), .CI(n1365), .CO(n708), .S(n709) );
  FADDX1 U421 ( .A(n1230), .B(n1418), .CI(n1250), .CO(n710), .S(n711) );
  FADDX1 U422 ( .A(n1193), .B(n1446), .CI(n1211), .CO(n712), .S(n713) );
  FADDX1 U423 ( .A(n1505), .B(n1340), .CI(n1475), .CO(n714), .S(n715) );
  FADDX1 U424 ( .A(n1160), .B(n1271), .CI(n1176), .CO(n716), .S(n717) );
  FADDX1 U425 ( .A(n1536), .B(n1316), .CI(n1145), .CO(n718), .S(n719) );
  HADDX1 U426 ( .A0(n1131), .B0(n1118), .C1(n720), .SO(n721) );
  FADDX1 U427 ( .A(n758), .B(n727), .CI(n725), .CO(n722), .S(n723) );
  FADDX1 U428 ( .A(n729), .B(n762), .CI(n760), .CO(n724), .S(n725) );
  FADDX1 U429 ( .A(n764), .B(n733), .CI(n731), .CO(n726), .S(n727) );
  FADDX1 U430 ( .A(n735), .B(n739), .CI(n766), .CO(n728), .S(n729) );
  FADDX1 U431 ( .A(n768), .B(n741), .CI(n737), .CO(n730), .S(n731) );
  FADDX1 U432 ( .A(n772), .B(n774), .CI(n770), .CO(n732), .S(n733) );
  FADDX1 U433 ( .A(n753), .B(n745), .CI(n743), .CO(n734), .S(n735) );
  FADDX1 U434 ( .A(n751), .B(n782), .CI(n747), .CO(n736), .S(n737) );
  FADDX1 U435 ( .A(n784), .B(n780), .CI(n749), .CO(n738), .S(n739) );
  FADDX1 U436 ( .A(n778), .B(n786), .CI(n776), .CO(n740), .S(n741) );
  FADDX1 U437 ( .A(n1366), .B(n1392), .CI(n755), .CO(n742), .S(n743) );
  FADDX1 U438 ( .A(n1251), .B(n1419), .CI(n1341), .CO(n744), .S(n745) );
  FADDX1 U439 ( .A(n1212), .B(n1447), .CI(n1231), .CO(n746), .S(n747) );
  FADDX1 U440 ( .A(n1476), .B(n1294), .CI(n1194), .CO(n748), .S(n749) );
  FADDX1 U441 ( .A(n1177), .B(n1272), .CI(n1506), .CO(n750), .S(n751) );
  FADDX1 U442 ( .A(n1537), .B(n1317), .CI(n1161), .CO(n752), .S(n753) );
  HADDX1 U443 ( .A0(n1146), .B0(n1132), .C1(n754), .SO(n755) );
  FADDX1 U444 ( .A(n790), .B(n761), .CI(n759), .CO(n756), .S(n757) );
  FADDX1 U445 ( .A(n763), .B(n765), .CI(n792), .CO(n758), .S(n759) );
  FADDX1 U446 ( .A(n796), .B(n767), .CI(n794), .CO(n760), .S(n761) );
  FADDX1 U447 ( .A(n769), .B(n773), .CI(n798), .CO(n762), .S(n763) );
  FADDX1 U448 ( .A(n800), .B(n802), .CI(n771), .CO(n764), .S(n765) );
  FADDX1 U449 ( .A(n775), .B(n785), .CI(n804), .CO(n766), .S(n767) );
  FADDX1 U450 ( .A(n781), .B(n810), .CI(n779), .CO(n768), .S(n769) );
  FADDX1 U451 ( .A(n812), .B(n806), .CI(n783), .CO(n770), .S(n771) );
  FADDX1 U452 ( .A(n814), .B(n808), .CI(n777), .CO(n772), .S(n773) );
  FADDX1 U453 ( .A(n787), .B(n1232), .CI(n816), .CO(n774), .S(n775) );
  FADDX1 U454 ( .A(n1318), .B(n1367), .CI(n1295), .CO(n776), .S(n777) );
  FADDX1 U455 ( .A(n1195), .B(n1393), .CI(n1213), .CO(n778), .S(n779) );
  FADDX1 U456 ( .A(n1178), .B(n1252), .CI(n1420), .CO(n780), .S(n781) );
  FADDX1 U457 ( .A(n1477), .B(n1273), .CI(n1448), .CO(n782), .S(n783) );
  FADDX1 U458 ( .A(n1538), .B(n1342), .CI(n1507), .CO(n784), .S(n785) );
  HADDX1 U459 ( .A0(n1162), .B0(n1147), .C1(n786), .SO(n787) );
  FADDX1 U460 ( .A(n820), .B(n793), .CI(n791), .CO(n788), .S(n789) );
  FADDX1 U461 ( .A(n795), .B(n797), .CI(n822), .CO(n790), .S(n791) );
  FADDX1 U462 ( .A(n826), .B(n799), .CI(n824), .CO(n792), .S(n793) );
  FADDX1 U463 ( .A(n803), .B(n828), .CI(n801), .CO(n794), .S(n795) );
  FADDX1 U464 ( .A(n832), .B(n805), .CI(n830), .CO(n796), .S(n797) );
  FADDX1 U465 ( .A(n815), .B(n807), .CI(n834), .CO(n798), .S(n799) );
  FADDX1 U466 ( .A(n813), .B(n838), .CI(n809), .CO(n800), .S(n801) );
  FADDX1 U467 ( .A(n840), .B(n836), .CI(n811), .CO(n802), .S(n803) );
  FADDX1 U468 ( .A(n844), .B(n817), .CI(n842), .CO(n804), .S(n805) );
  FADDX1 U469 ( .A(n1394), .B(n1274), .CI(n1319), .CO(n806), .S(n807) );
  FADDX1 U470 ( .A(n1233), .B(n1421), .CI(n1253), .CO(n808), .S(n809) );
  FADDX1 U471 ( .A(n1478), .B(n1296), .CI(n1449), .CO(n810), .S(n811) );
  FADDX1 U472 ( .A(n1539), .B(n1368), .CI(n1508), .CO(n812), .S(n813) );
  FADDX1 U473 ( .A(n1196), .B(n1343), .CI(n1214), .CO(n814), .S(n815) );
  HADDX1 U474 ( .A0(n1179), .B0(n1163), .C1(n816), .SO(n817) );
  FADDX1 U475 ( .A(n848), .B(n823), .CI(n821), .CO(n818), .S(n819) );
  FADDX1 U476 ( .A(n825), .B(n852), .CI(n850), .CO(n820), .S(n821) );
  FADDX1 U477 ( .A(n854), .B(n829), .CI(n827), .CO(n822), .S(n823) );
  FADDX1 U478 ( .A(n833), .B(n856), .CI(n831), .CO(n824), .S(n825) );
  FADDX1 U479 ( .A(n860), .B(n835), .CI(n858), .CO(n826), .S(n827) );
  FADDX1 U480 ( .A(n839), .B(n841), .CI(n837), .CO(n828), .S(n829) );
  FADDX1 U481 ( .A(n868), .B(n866), .CI(n843), .CO(n830), .S(n831) );
  FADDX1 U482 ( .A(n864), .B(n870), .CI(n862), .CO(n832), .S(n833) );
  FADDX1 U483 ( .A(n1395), .B(n1344), .CI(n845), .CO(n834), .S(n835) );
  FADDX1 U484 ( .A(n1275), .B(n1422), .CI(n1320), .CO(n836), .S(n837) );
  FADDX1 U485 ( .A(n1215), .B(n1254), .CI(n1234), .CO(n838), .S(n839) );
  FADDX1 U486 ( .A(n1479), .B(n1297), .CI(n1450), .CO(n840), .S(n841) );
  FADDX1 U487 ( .A(n1540), .B(n1369), .CI(n1509), .CO(n842), .S(n843) );
  HADDX1 U488 ( .A0(n1197), .B0(n1180), .C1(n844), .SO(n845) );
  FADDX1 U489 ( .A(n874), .B(n851), .CI(n849), .CO(n846), .S(n847) );
  FADDX1 U490 ( .A(n853), .B(n878), .CI(n876), .CO(n848), .S(n849) );
  FADDX1 U491 ( .A(n859), .B(n857), .CI(n855), .CO(n850), .S(n851) );
  FADDX1 U492 ( .A(n882), .B(n884), .CI(n880), .CO(n852), .S(n853) );
  FADDX1 U493 ( .A(n865), .B(n867), .CI(n861), .CO(n854), .S(n855) );
  FADDX1 U494 ( .A(n890), .B(n892), .CI(n869), .CO(n856), .S(n857) );
  FADDX1 U495 ( .A(n886), .B(n888), .CI(n863), .CO(n858), .S(n859) );
  FADDX1 U496 ( .A(n871), .B(n1451), .CI(n894), .CO(n860), .S(n861) );
  FADDX1 U497 ( .A(n1321), .B(n1480), .CI(n1423), .CO(n862), .S(n863) );
  FADDX1 U498 ( .A(n1510), .B(n1345), .CI(n1298), .CO(n864), .S(n865) );
  FADDX1 U499 ( .A(n1276), .B(n1396), .CI(n1541), .CO(n866), .S(n867) );
  FADDX1 U500 ( .A(n1235), .B(n1370), .CI(n1255), .CO(n868), .S(n869) );
  HADDX1 U501 ( .A0(n1216), .B0(n1198), .C1(n870), .SO(n871) );
  FADDX1 U502 ( .A(n898), .B(n877), .CI(n875), .CO(n872), .S(n873) );
  FADDX1 U503 ( .A(n879), .B(n902), .CI(n900), .CO(n874), .S(n875) );
  FADDX1 U504 ( .A(n883), .B(n904), .CI(n881), .CO(n876), .S(n877) );
  FADDX1 U505 ( .A(n885), .B(n908), .CI(n906), .CO(n878), .S(n879) );
  FADDX1 U506 ( .A(n891), .B(n887), .CI(n889), .CO(n880), .S(n881) );
  FADDX1 U507 ( .A(n910), .B(n912), .CI(n893), .CO(n882), .S(n883) );
  FADDX1 U508 ( .A(n916), .B(n895), .CI(n914), .CO(n884), .S(n885) );
  FADDX1 U509 ( .A(n1371), .B(n1452), .CI(n1424), .CO(n886), .S(n887) );
  FADDX1 U510 ( .A(n1299), .B(n1481), .CI(n1346), .CO(n888), .S(n889) );
  FADDX1 U511 ( .A(n1256), .B(n1322), .CI(n1277), .CO(n890), .S(n891) );
  FADDX1 U512 ( .A(n1542), .B(n1397), .CI(n1511), .CO(n892), .S(n893) );
  HADDX1 U513 ( .A0(n1236), .B0(n1217), .C1(n894), .SO(n895) );
  FADDX1 U514 ( .A(n920), .B(n901), .CI(n899), .CO(n896), .S(n897) );
  FADDX1 U515 ( .A(n903), .B(n905), .CI(n922), .CO(n898), .S(n899) );
  FADDX1 U516 ( .A(n907), .B(n926), .CI(n924), .CO(n900), .S(n901) );
  FADDX1 U517 ( .A(n909), .B(n913), .CI(n928), .CO(n902), .S(n903) );
  FADDX1 U518 ( .A(n911), .B(n930), .CI(n915), .CO(n904), .S(n905) );
  FADDX1 U519 ( .A(n934), .B(n936), .CI(n932), .CO(n906), .S(n907) );
  FADDX1 U520 ( .A(n1425), .B(n1453), .CI(n917), .CO(n908), .S(n909) );
  FADDX1 U521 ( .A(n1323), .B(n1482), .CI(n1347), .CO(n910), .S(n911) );
  FADDX1 U522 ( .A(n1543), .B(n1372), .CI(n1512), .CO(n912), .S(n913) );
  FADDX1 U523 ( .A(n1278), .B(n1398), .CI(n1300), .CO(n914), .S(n915) );
  HADDX1 U524 ( .A0(n1257), .B0(n1237), .C1(n916), .SO(n917) );
  FADDX1 U525 ( .A(n940), .B(n923), .CI(n921), .CO(n918), .S(n919) );
  FADDX1 U526 ( .A(n925), .B(n927), .CI(n942), .CO(n920), .S(n921) );
  FADDX1 U527 ( .A(n946), .B(n929), .CI(n944), .CO(n922), .S(n923) );
  FADDX1 U528 ( .A(n931), .B(n950), .CI(n935), .CO(n924), .S(n925) );
  FADDX1 U529 ( .A(n948), .B(n952), .CI(n933), .CO(n926), .S(n927) );
  FADDX1 U530 ( .A(n937), .B(n1454), .CI(n954), .CO(n928), .S(n929) );
  FADDX1 U531 ( .A(n1373), .B(n1483), .CI(n1426), .CO(n930), .S(n931) );
  FADDX1 U532 ( .A(n1301), .B(n1348), .CI(n1324), .CO(n932), .S(n933) );
  FADDX1 U533 ( .A(n1544), .B(n1399), .CI(n1513), .CO(n934), .S(n935) );
  HADDX1 U534 ( .A0(n1279), .B0(n1258), .C1(n936), .SO(n937) );
  FADDX1 U535 ( .A(n958), .B(n943), .CI(n941), .CO(n938), .S(n939) );
  FADDX1 U536 ( .A(n945), .B(n962), .CI(n960), .CO(n940), .S(n941) );
  FADDX1 U537 ( .A(n964), .B(n951), .CI(n947), .CO(n942), .S(n943) );
  FADDX1 U538 ( .A(n949), .B(n966), .CI(n953), .CO(n944), .S(n945) );
  FADDX1 U539 ( .A(n970), .B(n955), .CI(n968), .CO(n946), .S(n947) );
  FADDX1 U540 ( .A(n1400), .B(n1514), .CI(n1484), .CO(n948), .S(n949) );
  FADDX1 U541 ( .A(n1545), .B(n1455), .CI(n1374), .CO(n950), .S(n951) );
  FADDX1 U542 ( .A(n1325), .B(n1427), .CI(n1349), .CO(n952), .S(n953) );
  HADDX1 U543 ( .A0(n1302), .B0(n1280), .C1(n954), .SO(n955) );
  FADDX1 U544 ( .A(n974), .B(n961), .CI(n959), .CO(n956), .S(n957) );
  FADDX1 U545 ( .A(n976), .B(n978), .CI(n963), .CO(n958), .S(n959) );
  FADDX1 U546 ( .A(n969), .B(n967), .CI(n965), .CO(n960), .S(n961) );
  FADDX1 U547 ( .A(n982), .B(n984), .CI(n980), .CO(n962), .S(n963) );
  FADDX1 U548 ( .A(n1456), .B(n1485), .CI(n971), .CO(n964), .S(n965) );
  FADDX1 U549 ( .A(n1350), .B(n1375), .CI(n1401), .CO(n966), .S(n967) );
  FADDX1 U550 ( .A(n1546), .B(n1428), .CI(n1515), .CO(n968), .S(n969) );
  HADDX1 U551 ( .A0(n1326), .B0(n1303), .C1(n970), .SO(n971) );
  FADDX1 U552 ( .A(n988), .B(n977), .CI(n975), .CO(n972), .S(n973) );
  FADDX1 U553 ( .A(n979), .B(n981), .CI(n990), .CO(n974), .S(n975) );
  FADDX1 U554 ( .A(n992), .B(n994), .CI(n983), .CO(n976), .S(n977) );
  FADDX1 U555 ( .A(n985), .B(n1486), .CI(n996), .CO(n978), .S(n979) );
  FADDX1 U556 ( .A(n1516), .B(n1429), .CI(n1402), .CO(n980), .S(n981) );
  FADDX1 U557 ( .A(n1376), .B(n1457), .CI(n1547), .CO(n982), .S(n983) );
  HADDX1 U558 ( .A0(n1351), .B0(n1327), .C1(n984), .SO(n985) );
  FADDX1 U559 ( .A(n1000), .B(n991), .CI(n989), .CO(n986), .S(n987) );
  FADDX1 U560 ( .A(n995), .B(n993), .CI(n1002), .CO(n988), .S(n989) );
  FADDX1 U561 ( .A(n1006), .B(n997), .CI(n1004), .CO(n990), .S(n991) );
  FADDX1 U562 ( .A(n1403), .B(n1487), .CI(n1430), .CO(n992), .S(n993) );
  FADDX1 U563 ( .A(n1548), .B(n1458), .CI(n1517), .CO(n994), .S(n995) );
  HADDX1 U564 ( .A0(n1377), .B0(n1352), .C1(n996), .SO(n997) );
  FADDX1 U565 ( .A(n1010), .B(n1003), .CI(n1001), .CO(n998), .S(n999) );
  FADDX1 U566 ( .A(n1012), .B(n1014), .CI(n1005), .CO(n1000), .S(n1001) );
  FADDX1 U567 ( .A(n1459), .B(n1518), .CI(n1007), .CO(n1002), .S(n1003) );
  FADDX1 U568 ( .A(n1431), .B(n1488), .CI(n1549), .CO(n1004), .S(n1005) );
  HADDX1 U569 ( .A0(n1404), .B0(n1378), .C1(n1006), .SO(n1007) );
  FADDX1 U570 ( .A(n1013), .B(n1018), .CI(n1011), .CO(n1008), .S(n1009) );
  FADDX1 U571 ( .A(n1015), .B(n1550), .CI(n1020), .CO(n1010), .S(n1011) );
  FADDX1 U572 ( .A(n1460), .B(n1489), .CI(n1519), .CO(n1012), .S(n1013) );
  HADDX1 U573 ( .A0(n1432), .B0(n1405), .C1(n1014), .SO(n1015) );
  FADDX1 U574 ( .A(n1024), .B(n1021), .CI(n1019), .CO(n1016), .S(n1017) );
  FADDX1 U575 ( .A(n1490), .B(n1551), .CI(n1520), .CO(n1018), .S(n1019) );
  HADDX1 U576 ( .A0(n1461), .B0(n1433), .C1(n1020), .SO(n1021) );
  FADDX1 U577 ( .A(n1521), .B(n1552), .CI(n1025), .CO(n1022), .S(n1023) );
  HADDX1 U578 ( .A0(n1491), .B0(n1462), .C1(n1024), .SO(n1025) );
  HADDX1 U579 ( .A0(n1553), .B0(n1522), .C1(n1026), .SO(n1027) );
  NOR2X0 U580 ( .IN1(n50), .IN2(n48), .QN(n1028) );
  NOR2X0 U581 ( .IN1(n1578), .IN2(n47), .QN(n1029) );
  NOR2X0 U582 ( .IN1(n50), .IN2(n47), .QN(n1030) );
  NOR2X0 U583 ( .IN1(n1577), .IN2(n46), .QN(n1031) );
  NOR2X0 U584 ( .IN1(n1578), .IN2(n46), .QN(n1032) );
  NOR2X0 U585 ( .IN1(n50), .IN2(n46), .QN(n1033) );
  NOR2X0 U586 ( .IN1(n1576), .IN2(n45), .QN(n1034) );
  NOR2X0 U587 ( .IN1(n1577), .IN2(n45), .QN(n1035) );
  NOR2X0 U588 ( .IN1(n1578), .IN2(n45), .QN(n1036) );
  NOR2X0 U589 ( .IN1(n50), .IN2(n45), .QN(n1037) );
  NOR2X0 U590 ( .IN1(n1575), .IN2(n1580), .QN(n1038) );
  NOR2X0 U591 ( .IN1(n1576), .IN2(n1580), .QN(n1039) );
  NOR2X0 U592 ( .IN1(n1577), .IN2(n1580), .QN(n1040) );
  NOR2X0 U593 ( .IN1(n1578), .IN2(n1580), .QN(n1041) );
  NOR2X0 U594 ( .IN1(n50), .IN2(n1580), .QN(n1042) );
  NOR2X0 U595 ( .IN1(n1574), .IN2(n1581), .QN(n1043) );
  NOR2X0 U596 ( .IN1(n1575), .IN2(n1581), .QN(n1044) );
  NOR2X0 U597 ( .IN1(n1576), .IN2(n1581), .QN(n1045) );
  NOR2X0 U598 ( .IN1(n1577), .IN2(n1581), .QN(n1046) );
  NOR2X0 U599 ( .IN1(n1578), .IN2(n1581), .QN(n1047) );
  NOR2X0 U600 ( .IN1(n50), .IN2(n1581), .QN(n1048) );
  NOR2X0 U601 ( .IN1(n62), .IN2(n1582), .QN(n1049) );
  NOR2X0 U602 ( .IN1(n1574), .IN2(n1582), .QN(n1050) );
  NOR2X0 U603 ( .IN1(n1575), .IN2(n1582), .QN(n1051) );
  NOR2X0 U604 ( .IN1(n1576), .IN2(n1582), .QN(n1052) );
  NOR2X0 U605 ( .IN1(n1577), .IN2(n1582), .QN(n1053) );
  NOR2X0 U606 ( .IN1(n1578), .IN2(n1582), .QN(n1054) );
  NOR2X0 U607 ( .IN1(n50), .IN2(n1582), .QN(n1055) );
  NOR2X0 U608 ( .IN1(n64), .IN2(n1583), .QN(n1056) );
  NOR2X0 U609 ( .IN1(n62), .IN2(n1583), .QN(n1057) );
  NOR2X0 U610 ( .IN1(n1574), .IN2(n1583), .QN(n1058) );
  NOR2X0 U611 ( .IN1(n1575), .IN2(n1583), .QN(n1059) );
  NOR2X0 U612 ( .IN1(n1576), .IN2(n1583), .QN(n1060) );
  NOR2X0 U613 ( .IN1(n1577), .IN2(n1583), .QN(n1061) );
  NOR2X0 U614 ( .IN1(n1578), .IN2(n1583), .QN(n1062) );
  NOR2X0 U615 ( .IN1(n50), .IN2(n1583), .QN(n1063) );
  NOR2X0 U616 ( .IN1(n1571), .IN2(n1584), .QN(n1064) );
  NOR2X0 U617 ( .IN1(n64), .IN2(n1584), .QN(n1065) );
  NOR2X0 U618 ( .IN1(n62), .IN2(n1584), .QN(n1066) );
  NOR2X0 U619 ( .IN1(n1574), .IN2(n1584), .QN(n1067) );
  NOR2X0 U620 ( .IN1(n1575), .IN2(n1584), .QN(n1068) );
  NOR2X0 U621 ( .IN1(n1576), .IN2(n1584), .QN(n1069) );
  NOR2X0 U622 ( .IN1(n1577), .IN2(n1584), .QN(n1070) );
  NOR2X0 U623 ( .IN1(n1578), .IN2(n1584), .QN(n1071) );
  NOR2X0 U624 ( .IN1(n50), .IN2(n1584), .QN(n1072) );
  NOR2X0 U625 ( .IN1(n1570), .IN2(n1585), .QN(n1073) );
  NOR2X0 U626 ( .IN1(n1571), .IN2(n1585), .QN(n1074) );
  NOR2X0 U627 ( .IN1(n64), .IN2(n1585), .QN(n1075) );
  NOR2X0 U628 ( .IN1(n62), .IN2(n1585), .QN(n1076) );
  NOR2X0 U629 ( .IN1(n1574), .IN2(n1585), .QN(n1077) );
  NOR2X0 U630 ( .IN1(n1575), .IN2(n1585), .QN(n1078) );
  NOR2X0 U631 ( .IN1(n1576), .IN2(n1585), .QN(n1079) );
  NOR2X0 U632 ( .IN1(n1577), .IN2(n1585), .QN(n1080) );
  NOR2X0 U633 ( .IN1(n1578), .IN2(n1585), .QN(n1081) );
  NOR2X0 U634 ( .IN1(n50), .IN2(n1585), .QN(n1082) );
  NOR2X0 U635 ( .IN1(n1569), .IN2(n1586), .QN(n1083) );
  NOR2X0 U636 ( .IN1(n1570), .IN2(n1586), .QN(n1084) );
  NOR2X0 U637 ( .IN1(n1571), .IN2(n1586), .QN(n1085) );
  NOR2X0 U638 ( .IN1(n64), .IN2(n1586), .QN(n1086) );
  NOR2X0 U639 ( .IN1(n62), .IN2(n1586), .QN(n1087) );
  NOR2X0 U640 ( .IN1(n1574), .IN2(n1586), .QN(n1088) );
  NOR2X0 U641 ( .IN1(n1575), .IN2(n1586), .QN(n1089) );
  NOR2X0 U642 ( .IN1(n1576), .IN2(n1586), .QN(n1090) );
  NOR2X0 U643 ( .IN1(n1577), .IN2(n1586), .QN(n1091) );
  NOR2X0 U644 ( .IN1(n1578), .IN2(n1586), .QN(n1092) );
  NOR2X0 U645 ( .IN1(n50), .IN2(n1586), .QN(n1093) );
  NOR2X0 U646 ( .IN1(n1568), .IN2(n1587), .QN(n1094) );
  NOR2X0 U647 ( .IN1(n1569), .IN2(n1587), .QN(n1095) );
  NOR2X0 U648 ( .IN1(n1570), .IN2(n1587), .QN(n1096) );
  NOR2X0 U649 ( .IN1(n1571), .IN2(n1587), .QN(n1097) );
  NOR2X0 U650 ( .IN1(n64), .IN2(n1587), .QN(n1098) );
  NOR2X0 U651 ( .IN1(n62), .IN2(n1587), .QN(n1099) );
  NOR2X0 U652 ( .IN1(n1574), .IN2(n1587), .QN(n1100) );
  NOR2X0 U653 ( .IN1(n1575), .IN2(n1587), .QN(n1101) );
  NOR2X0 U654 ( .IN1(n1576), .IN2(n1587), .QN(n1102) );
  NOR2X0 U655 ( .IN1(n1577), .IN2(n1587), .QN(n1103) );
  NOR2X0 U656 ( .IN1(n1578), .IN2(n1587), .QN(n1104) );
  NOR2X0 U657 ( .IN1(n50), .IN2(n1587), .QN(n1105) );
  NOR2X0 U658 ( .IN1(n74), .IN2(n1588), .QN(n1106) );
  NOR2X0 U659 ( .IN1(n1568), .IN2(n1588), .QN(n1107) );
  NOR2X0 U660 ( .IN1(n1569), .IN2(n1588), .QN(n1108) );
  NOR2X0 U661 ( .IN1(n1570), .IN2(n1588), .QN(n1109) );
  NOR2X0 U662 ( .IN1(n1571), .IN2(n1588), .QN(n1110) );
  NOR2X0 U663 ( .IN1(n64), .IN2(n1588), .QN(n1111) );
  NOR2X0 U664 ( .IN1(n62), .IN2(n1588), .QN(n1112) );
  NOR2X0 U665 ( .IN1(n1574), .IN2(n1588), .QN(n1113) );
  NOR2X0 U666 ( .IN1(n1575), .IN2(n1588), .QN(n1114) );
  NOR2X0 U667 ( .IN1(n1576), .IN2(n1588), .QN(n1115) );
  NOR2X0 U668 ( .IN1(n1577), .IN2(n1588), .QN(n1116) );
  NOR2X0 U669 ( .IN1(n1578), .IN2(n1588), .QN(n1117) );
  NOR2X0 U670 ( .IN1(n50), .IN2(n1588), .QN(n1118) );
  NOR2X0 U671 ( .IN1(n76), .IN2(n1589), .QN(n1119) );
  NOR2X0 U672 ( .IN1(n74), .IN2(n1589), .QN(n1120) );
  NOR2X0 U673 ( .IN1(n1568), .IN2(n1589), .QN(n1121) );
  NOR2X0 U674 ( .IN1(n1569), .IN2(n1589), .QN(n1122) );
  NOR2X0 U675 ( .IN1(n1570), .IN2(n1589), .QN(n1123) );
  NOR2X0 U676 ( .IN1(n1571), .IN2(n1589), .QN(n1124) );
  NOR2X0 U677 ( .IN1(n64), .IN2(n1589), .QN(n1125) );
  NOR2X0 U678 ( .IN1(n62), .IN2(n1589), .QN(n1126) );
  NOR2X0 U679 ( .IN1(n1574), .IN2(n1589), .QN(n1127) );
  NOR2X0 U680 ( .IN1(n1575), .IN2(n1589), .QN(n1128) );
  NOR2X0 U681 ( .IN1(n1576), .IN2(n1589), .QN(n1129) );
  NOR2X0 U682 ( .IN1(n1577), .IN2(n1589), .QN(n1130) );
  NOR2X0 U683 ( .IN1(n1578), .IN2(n1589), .QN(n1131) );
  NOR2X0 U684 ( .IN1(n50), .IN2(n1589), .QN(n1132) );
  NOR2X0 U685 ( .IN1(n78), .IN2(n1590), .QN(n1133) );
  NOR2X0 U686 ( .IN1(n76), .IN2(n1590), .QN(n1134) );
  NOR2X0 U687 ( .IN1(n74), .IN2(n1590), .QN(n1135) );
  NOR2X0 U688 ( .IN1(n1568), .IN2(n1590), .QN(n1136) );
  NOR2X0 U689 ( .IN1(n1569), .IN2(n1590), .QN(n1137) );
  NOR2X0 U690 ( .IN1(n1570), .IN2(n1590), .QN(n1138) );
  NOR2X0 U691 ( .IN1(n1571), .IN2(n1590), .QN(n1139) );
  NOR2X0 U692 ( .IN1(n64), .IN2(n1590), .QN(n1140) );
  NOR2X0 U693 ( .IN1(n62), .IN2(n1590), .QN(n1141) );
  NOR2X0 U694 ( .IN1(n1574), .IN2(n1590), .QN(n1142) );
  NOR2X0 U695 ( .IN1(n1575), .IN2(n1590), .QN(n1143) );
  NOR2X0 U696 ( .IN1(n1576), .IN2(n1590), .QN(n1144) );
  NOR2X0 U697 ( .IN1(n1577), .IN2(n1590), .QN(n1145) );
  NOR2X0 U698 ( .IN1(n1578), .IN2(n1590), .QN(n1146) );
  NOR2X0 U699 ( .IN1(n50), .IN2(n1590), .QN(n1147) );
  NOR2X0 U700 ( .IN1(n80), .IN2(n1591), .QN(n1148) );
  NOR2X0 U701 ( .IN1(n78), .IN2(n1591), .QN(n1149) );
  NOR2X0 U702 ( .IN1(n76), .IN2(n1591), .QN(n1150) );
  NOR2X0 U703 ( .IN1(n74), .IN2(n1591), .QN(n1151) );
  NOR2X0 U704 ( .IN1(n1568), .IN2(n1591), .QN(n1152) );
  NOR2X0 U705 ( .IN1(n1569), .IN2(n1591), .QN(n1153) );
  NOR2X0 U706 ( .IN1(n1570), .IN2(n1591), .QN(n1154) );
  NOR2X0 U707 ( .IN1(n1571), .IN2(n1591), .QN(n1155) );
  NOR2X0 U708 ( .IN1(n64), .IN2(n1591), .QN(n1156) );
  NOR2X0 U709 ( .IN1(n62), .IN2(n1591), .QN(n1157) );
  NOR2X0 U710 ( .IN1(n1574), .IN2(n1591), .QN(n1158) );
  NOR2X0 U711 ( .IN1(n1575), .IN2(n1591), .QN(n1159) );
  NOR2X0 U712 ( .IN1(n1576), .IN2(n1591), .QN(n1160) );
  NOR2X0 U713 ( .IN1(n1577), .IN2(n1591), .QN(n1161) );
  NOR2X0 U714 ( .IN1(n1578), .IN2(n1591), .QN(n1162) );
  NOR2X0 U715 ( .IN1(n50), .IN2(n1591), .QN(n1163) );
  NOR2X0 U716 ( .IN1(n1566), .IN2(n32), .QN(n1164) );
  NOR2X0 U717 ( .IN1(n80), .IN2(n32), .QN(n1165) );
  NOR2X0 U718 ( .IN1(n78), .IN2(n32), .QN(n1166) );
  NOR2X0 U719 ( .IN1(n76), .IN2(n32), .QN(n1167) );
  NOR2X0 U720 ( .IN1(n74), .IN2(n32), .QN(n1168) );
  NOR2X0 U721 ( .IN1(n1568), .IN2(n32), .QN(n1169) );
  NOR2X0 U722 ( .IN1(n69), .IN2(n32), .QN(n1170) );
  NOR2X0 U723 ( .IN1(n67), .IN2(n32), .QN(n1171) );
  NOR2X0 U724 ( .IN1(n65), .IN2(n32), .QN(n1172) );
  NOR2X0 U725 ( .IN1(n1572), .IN2(n32), .QN(n1173) );
  NOR2X0 U726 ( .IN1(n62), .IN2(n32), .QN(n1174) );
  NOR2X0 U727 ( .IN1(n59), .IN2(n32), .QN(n1175) );
  NOR2X0 U728 ( .IN1(n57), .IN2(n32), .QN(n1176) );
  NOR2X0 U729 ( .IN1(n55), .IN2(n32), .QN(n1177) );
  NOR2X0 U730 ( .IN1(n53), .IN2(n32), .QN(n1178) );
  NOR2X0 U731 ( .IN1(n51), .IN2(n32), .QN(n1179) );
  NOR2X0 U732 ( .IN1(n50), .IN2(n32), .QN(n1180) );
  NOR2X0 U733 ( .IN1(n1565), .IN2(n30), .QN(n1181) );
  NOR2X0 U734 ( .IN1(n1566), .IN2(n30), .QN(n1182) );
  NOR2X0 U735 ( .IN1(n80), .IN2(n30), .QN(n1183) );
  NOR2X0 U736 ( .IN1(n78), .IN2(n30), .QN(n1184) );
  NOR2X0 U737 ( .IN1(n76), .IN2(n30), .QN(n1185) );
  NOR2X0 U738 ( .IN1(n1567), .IN2(n30), .QN(n1186) );
  NOR2X0 U739 ( .IN1(n1568), .IN2(n30), .QN(n1187) );
  NOR2X0 U740 ( .IN1(n69), .IN2(n30), .QN(n1188) );
  NOR2X0 U741 ( .IN1(n67), .IN2(n30), .QN(n1189) );
  NOR2X0 U742 ( .IN1(n65), .IN2(n30), .QN(n1190) );
  NOR2X0 U743 ( .IN1(n64), .IN2(n30), .QN(n1191) );
  NOR2X0 U744 ( .IN1(n1573), .IN2(n30), .QN(n1192) );
  NOR2X0 U745 ( .IN1(n59), .IN2(n30), .QN(n1193) );
  NOR2X0 U746 ( .IN1(n57), .IN2(n30), .QN(n1194) );
  NOR2X0 U747 ( .IN1(n55), .IN2(n30), .QN(n1195) );
  NOR2X0 U748 ( .IN1(n53), .IN2(n30), .QN(n1196) );
  NOR2X0 U749 ( .IN1(n51), .IN2(n30), .QN(n1197) );
  NOR2X0 U750 ( .IN1(n1579), .IN2(n30), .QN(n1198) );
  NOR2X0 U751 ( .IN1(n1564), .IN2(n28), .QN(n1199) );
  NOR2X0 U752 ( .IN1(n1565), .IN2(n28), .QN(n1200) );
  NOR2X0 U753 ( .IN1(n1566), .IN2(n28), .QN(n1201) );
  NOR2X0 U754 ( .IN1(n80), .IN2(n28), .QN(n1202) );
  NOR2X0 U755 ( .IN1(n78), .IN2(n28), .QN(n1203) );
  NOR2X0 U756 ( .IN1(n76), .IN2(n28), .QN(n1204) );
  NOR2X0 U757 ( .IN1(n74), .IN2(n28), .QN(n1205) );
  NOR2X0 U758 ( .IN1(n1568), .IN2(n28), .QN(n1206) );
  NOR2X0 U759 ( .IN1(n69), .IN2(n28), .QN(n1207) );
  NOR2X0 U760 ( .IN1(n67), .IN2(n28), .QN(n1208) );
  NOR2X0 U761 ( .IN1(n65), .IN2(n28), .QN(n1209) );
  NOR2X0 U762 ( .IN1(n1572), .IN2(n28), .QN(n1210) );
  NOR2X0 U763 ( .IN1(n62), .IN2(n28), .QN(n1211) );
  NOR2X0 U764 ( .IN1(n59), .IN2(n28), .QN(n1212) );
  NOR2X0 U765 ( .IN1(n57), .IN2(n28), .QN(n1213) );
  NOR2X0 U766 ( .IN1(n55), .IN2(n28), .QN(n1214) );
  NOR2X0 U767 ( .IN1(n53), .IN2(n28), .QN(n1215) );
  NOR2X0 U768 ( .IN1(n51), .IN2(n28), .QN(n1216) );
  NOR2X0 U769 ( .IN1(n1579), .IN2(n28), .QN(n1217) );
  NOR2X0 U770 ( .IN1(n1563), .IN2(n1592), .QN(n1218) );
  NOR2X0 U771 ( .IN1(n1564), .IN2(n1592), .QN(n1219) );
  NOR2X0 U772 ( .IN1(n1565), .IN2(n1592), .QN(n1220) );
  NOR2X0 U773 ( .IN1(n1566), .IN2(n1592), .QN(n1221) );
  NOR2X0 U774 ( .IN1(n80), .IN2(n1592), .QN(n1222) );
  NOR2X0 U775 ( .IN1(n78), .IN2(n1592), .QN(n1223) );
  NOR2X0 U776 ( .IN1(n76), .IN2(n1592), .QN(n1224) );
  NOR2X0 U777 ( .IN1(n1567), .IN2(n1592), .QN(n1225) );
  NOR2X0 U778 ( .IN1(n1568), .IN2(n1592), .QN(n1226) );
  NOR2X0 U779 ( .IN1(n69), .IN2(n1592), .QN(n1227) );
  NOR2X0 U780 ( .IN1(n67), .IN2(n1592), .QN(n1228) );
  NOR2X0 U781 ( .IN1(n65), .IN2(n1592), .QN(n1229) );
  NOR2X0 U782 ( .IN1(n64), .IN2(n1592), .QN(n1230) );
  NOR2X0 U783 ( .IN1(n1573), .IN2(n1592), .QN(n1231) );
  NOR2X0 U784 ( .IN1(n59), .IN2(n1592), .QN(n1232) );
  NOR2X0 U785 ( .IN1(n57), .IN2(n1592), .QN(n1233) );
  NOR2X0 U786 ( .IN1(n55), .IN2(n1592), .QN(n1234) );
  NOR2X0 U787 ( .IN1(n53), .IN2(n1592), .QN(n1235) );
  NOR2X0 U788 ( .IN1(n51), .IN2(n1592), .QN(n1236) );
  NOR2X0 U789 ( .IN1(n1579), .IN2(n1592), .QN(n1237) );
  NOR2X0 U790 ( .IN1(n1562), .IN2(n24), .QN(n1238) );
  NOR2X0 U791 ( .IN1(n1563), .IN2(n24), .QN(n1239) );
  NOR2X0 U792 ( .IN1(n1564), .IN2(n24), .QN(n1240) );
  NOR2X0 U793 ( .IN1(n1565), .IN2(n24), .QN(n1241) );
  NOR2X0 U794 ( .IN1(n1566), .IN2(n24), .QN(n1242) );
  NOR2X0 U795 ( .IN1(n80), .IN2(n1593), .QN(n1243) );
  NOR2X0 U796 ( .IN1(n78), .IN2(n24), .QN(n1244) );
  NOR2X0 U797 ( .IN1(n76), .IN2(n1593), .QN(n1245) );
  NOR2X0 U798 ( .IN1(n1567), .IN2(n24), .QN(n1246) );
  NOR2X0 U799 ( .IN1(n1568), .IN2(n1593), .QN(n1247) );
  NOR2X0 U800 ( .IN1(n69), .IN2(n1593), .QN(n1248) );
  NOR2X0 U801 ( .IN1(n67), .IN2(n24), .QN(n1249) );
  NOR2X0 U802 ( .IN1(n65), .IN2(n1593), .QN(n1250) );
  NOR2X0 U803 ( .IN1(n1572), .IN2(n24), .QN(n1251) );
  NOR2X0 U804 ( .IN1(n62), .IN2(n1593), .QN(n1252) );
  NOR2X0 U805 ( .IN1(n59), .IN2(n24), .QN(n1253) );
  NOR2X0 U806 ( .IN1(n57), .IN2(n1593), .QN(n1254) );
  NOR2X0 U807 ( .IN1(n55), .IN2(n24), .QN(n1255) );
  NOR2X0 U808 ( .IN1(n53), .IN2(n1593), .QN(n1256) );
  NOR2X0 U809 ( .IN1(n51), .IN2(n1593), .QN(n1257) );
  NOR2X0 U810 ( .IN1(n1579), .IN2(n1593), .QN(n1258) );
  NOR2X0 U811 ( .IN1(n1561), .IN2(n1594), .QN(n1259) );
  NOR2X0 U812 ( .IN1(n1562), .IN2(n1594), .QN(n1260) );
  NOR2X0 U813 ( .IN1(n1563), .IN2(n1594), .QN(n1261) );
  NOR2X0 U814 ( .IN1(n1564), .IN2(n1594), .QN(n1262) );
  NOR2X0 U815 ( .IN1(n1565), .IN2(n1594), .QN(n1263) );
  NOR2X0 U816 ( .IN1(n1566), .IN2(n1594), .QN(n1264) );
  NOR2X0 U817 ( .IN1(n80), .IN2(n21), .QN(n1265) );
  NOR2X0 U818 ( .IN1(n78), .IN2(n21), .QN(n1266) );
  NOR2X0 U819 ( .IN1(n76), .IN2(n21), .QN(n1267) );
  NOR2X0 U820 ( .IN1(n1567), .IN2(n21), .QN(n1268) );
  NOR2X0 U821 ( .IN1(n1568), .IN2(n21), .QN(n1269) );
  NOR2X0 U822 ( .IN1(n69), .IN2(n21), .QN(n1270) );
  NOR2X0 U823 ( .IN1(n67), .IN2(n21), .QN(n1271) );
  NOR2X0 U824 ( .IN1(n65), .IN2(n21), .QN(n1272) );
  NOR2X0 U825 ( .IN1(n64), .IN2(n21), .QN(n1273) );
  NOR2X0 U826 ( .IN1(n1573), .IN2(n21), .QN(n1274) );
  NOR2X0 U827 ( .IN1(n59), .IN2(n21), .QN(n1275) );
  NOR2X0 U828 ( .IN1(n57), .IN2(n21), .QN(n1276) );
  NOR2X0 U829 ( .IN1(n55), .IN2(n21), .QN(n1277) );
  NOR2X0 U830 ( .IN1(n53), .IN2(n21), .QN(n1278) );
  NOR2X0 U831 ( .IN1(n51), .IN2(n21), .QN(n1279) );
  NOR2X0 U832 ( .IN1(n1579), .IN2(n21), .QN(n1280) );
  NOR2X0 U833 ( .IN1(n1560), .IN2(n1595), .QN(n1281) );
  NOR2X0 U834 ( .IN1(n1561), .IN2(n1595), .QN(n1282) );
  NOR2X0 U835 ( .IN1(n1562), .IN2(n1595), .QN(n1283) );
  NOR2X0 U836 ( .IN1(n1563), .IN2(n1595), .QN(n1284) );
  NOR2X0 U837 ( .IN1(n1564), .IN2(n1595), .QN(n1285) );
  NOR2X0 U838 ( .IN1(n1565), .IN2(n1595), .QN(n1286) );
  NOR2X0 U839 ( .IN1(n1566), .IN2(n1595), .QN(n1287) );
  NOR2X0 U840 ( .IN1(n80), .IN2(n19), .QN(n1288) );
  NOR2X0 U841 ( .IN1(n78), .IN2(n19), .QN(n1289) );
  NOR2X0 U842 ( .IN1(n76), .IN2(n19), .QN(n1290) );
  NOR2X0 U843 ( .IN1(n74), .IN2(n19), .QN(n1291) );
  NOR2X0 U844 ( .IN1(n1568), .IN2(n19), .QN(n1292) );
  NOR2X0 U845 ( .IN1(n69), .IN2(n19), .QN(n1293) );
  NOR2X0 U846 ( .IN1(n67), .IN2(n19), .QN(n1294) );
  NOR2X0 U847 ( .IN1(n65), .IN2(n19), .QN(n1295) );
  NOR2X0 U848 ( .IN1(n1572), .IN2(n19), .QN(n1296) );
  NOR2X0 U849 ( .IN1(n62), .IN2(n19), .QN(n1297) );
  NOR2X0 U850 ( .IN1(n59), .IN2(n19), .QN(n1298) );
  NOR2X0 U851 ( .IN1(n57), .IN2(n19), .QN(n1299) );
  NOR2X0 U852 ( .IN1(n55), .IN2(n19), .QN(n1300) );
  NOR2X0 U853 ( .IN1(n53), .IN2(n19), .QN(n1301) );
  NOR2X0 U854 ( .IN1(n51), .IN2(n19), .QN(n1302) );
  NOR2X0 U855 ( .IN1(n1579), .IN2(n19), .QN(n1303) );
  NOR2X0 U856 ( .IN1(n1559), .IN2(n1596), .QN(n1304) );
  NOR2X0 U857 ( .IN1(n1560), .IN2(n1596), .QN(n1305) );
  NOR2X0 U858 ( .IN1(n1561), .IN2(n1596), .QN(n1306) );
  NOR2X0 U859 ( .IN1(n1562), .IN2(n1596), .QN(n1307) );
  NOR2X0 U860 ( .IN1(n1563), .IN2(n1596), .QN(n1308) );
  NOR2X0 U861 ( .IN1(n1564), .IN2(n1596), .QN(n1309) );
  NOR2X0 U862 ( .IN1(n1565), .IN2(n1596), .QN(n1310) );
  NOR2X0 U863 ( .IN1(n1566), .IN2(n1596), .QN(n1311) );
  NOR2X0 U864 ( .IN1(n80), .IN2(n17), .QN(n1312) );
  NOR2X0 U865 ( .IN1(n78), .IN2(n17), .QN(n1313) );
  NOR2X0 U866 ( .IN1(n76), .IN2(n17), .QN(n1314) );
  NOR2X0 U867 ( .IN1(n1567), .IN2(n17), .QN(n1315) );
  NOR2X0 U868 ( .IN1(n1568), .IN2(n17), .QN(n1316) );
  NOR2X0 U869 ( .IN1(n69), .IN2(n17), .QN(n1317) );
  NOR2X0 U870 ( .IN1(n67), .IN2(n17), .QN(n1318) );
  NOR2X0 U871 ( .IN1(n65), .IN2(n17), .QN(n1319) );
  NOR2X0 U872 ( .IN1(n64), .IN2(n17), .QN(n1320) );
  NOR2X0 U873 ( .IN1(n1573), .IN2(n17), .QN(n1321) );
  NOR2X0 U874 ( .IN1(n59), .IN2(n17), .QN(n1322) );
  NOR2X0 U875 ( .IN1(n57), .IN2(n17), .QN(n1323) );
  NOR2X0 U876 ( .IN1(n55), .IN2(n17), .QN(n1324) );
  NOR2X0 U877 ( .IN1(n53), .IN2(n17), .QN(n1325) );
  NOR2X0 U878 ( .IN1(n51), .IN2(n17), .QN(n1326) );
  NOR2X0 U879 ( .IN1(n1579), .IN2(n17), .QN(n1327) );
  NOR2X0 U880 ( .IN1(n1558), .IN2(n1597), .QN(n1328) );
  NOR2X0 U881 ( .IN1(n1559), .IN2(n1597), .QN(n1329) );
  NOR2X0 U882 ( .IN1(n1560), .IN2(n1597), .QN(n1330) );
  NOR2X0 U883 ( .IN1(n1561), .IN2(n1597), .QN(n1331) );
  NOR2X0 U884 ( .IN1(n1562), .IN2(n1597), .QN(n1332) );
  NOR2X0 U885 ( .IN1(n1563), .IN2(n1597), .QN(n1333) );
  NOR2X0 U886 ( .IN1(n1564), .IN2(n1597), .QN(n1334) );
  NOR2X0 U887 ( .IN1(n1565), .IN2(n1597), .QN(n1335) );
  NOR2X0 U888 ( .IN1(n1566), .IN2(n1597), .QN(n1336) );
  NOR2X0 U889 ( .IN1(n80), .IN2(n15), .QN(n1337) );
  NOR2X0 U890 ( .IN1(n78), .IN2(n15), .QN(n1338) );
  NOR2X0 U891 ( .IN1(n76), .IN2(n15), .QN(n1339) );
  NOR2X0 U892 ( .IN1(n74), .IN2(n15), .QN(n1340) );
  NOR2X0 U893 ( .IN1(n1568), .IN2(n15), .QN(n1341) );
  NOR2X0 U894 ( .IN1(n69), .IN2(n15), .QN(n1342) );
  NOR2X0 U895 ( .IN1(n67), .IN2(n15), .QN(n1343) );
  NOR2X0 U896 ( .IN1(n65), .IN2(n15), .QN(n1344) );
  NOR2X0 U897 ( .IN1(n1572), .IN2(n15), .QN(n1345) );
  NOR2X0 U898 ( .IN1(n1573), .IN2(n15), .QN(n1346) );
  NOR2X0 U899 ( .IN1(n59), .IN2(n15), .QN(n1347) );
  NOR2X0 U900 ( .IN1(n57), .IN2(n15), .QN(n1348) );
  NOR2X0 U901 ( .IN1(n55), .IN2(n15), .QN(n1349) );
  NOR2X0 U902 ( .IN1(n53), .IN2(n15), .QN(n1350) );
  NOR2X0 U903 ( .IN1(n51), .IN2(n15), .QN(n1351) );
  NOR2X0 U904 ( .IN1(n1579), .IN2(n15), .QN(n1352) );
  NOR2X0 U905 ( .IN1(n1557), .IN2(n1598), .QN(n1353) );
  NOR2X0 U906 ( .IN1(n1558), .IN2(n1598), .QN(n1354) );
  NOR2X0 U907 ( .IN1(n1559), .IN2(n1598), .QN(n1355) );
  NOR2X0 U908 ( .IN1(n1560), .IN2(n1598), .QN(n1356) );
  NOR2X0 U909 ( .IN1(n1561), .IN2(n1598), .QN(n1357) );
  NOR2X0 U910 ( .IN1(n1562), .IN2(n1598), .QN(n1358) );
  NOR2X0 U911 ( .IN1(n1563), .IN2(n1598), .QN(n1359) );
  NOR2X0 U912 ( .IN1(n1564), .IN2(n1598), .QN(n1360) );
  NOR2X0 U913 ( .IN1(n1565), .IN2(n1598), .QN(n1361) );
  NOR2X0 U914 ( .IN1(n1566), .IN2(n1598), .QN(n1362) );
  NOR2X0 U915 ( .IN1(n80), .IN2(n13), .QN(n1363) );
  NOR2X0 U916 ( .IN1(n78), .IN2(n13), .QN(n1364) );
  NOR2X0 U917 ( .IN1(n76), .IN2(n13), .QN(n1365) );
  NOR2X0 U918 ( .IN1(n1567), .IN2(n13), .QN(n1366) );
  NOR2X0 U919 ( .IN1(n1568), .IN2(n13), .QN(n1367) );
  NOR2X0 U920 ( .IN1(n69), .IN2(n13), .QN(n1368) );
  NOR2X0 U921 ( .IN1(n67), .IN2(n13), .QN(n1369) );
  NOR2X0 U922 ( .IN1(n65), .IN2(n13), .QN(n1370) );
  NOR2X0 U923 ( .IN1(n1572), .IN2(n13), .QN(n1371) );
  NOR2X0 U924 ( .IN1(n1573), .IN2(n13), .QN(n1372) );
  NOR2X0 U925 ( .IN1(n59), .IN2(n13), .QN(n1373) );
  NOR2X0 U926 ( .IN1(n57), .IN2(n13), .QN(n1374) );
  NOR2X0 U927 ( .IN1(n55), .IN2(n13), .QN(n1375) );
  NOR2X0 U928 ( .IN1(n53), .IN2(n13), .QN(n1376) );
  NOR2X0 U929 ( .IN1(n51), .IN2(n13), .QN(n1377) );
  NOR2X0 U930 ( .IN1(n1579), .IN2(n13), .QN(n1378) );
  NOR2X0 U931 ( .IN1(n1556), .IN2(n12), .QN(n1379) );
  NOR2X0 U932 ( .IN1(n1557), .IN2(n12), .QN(n1380) );
  NOR2X0 U933 ( .IN1(n1558), .IN2(n12), .QN(n1381) );
  NOR2X0 U934 ( .IN1(n1559), .IN2(n12), .QN(n1382) );
  NOR2X0 U935 ( .IN1(n1560), .IN2(n12), .QN(n1383) );
  NOR2X0 U936 ( .IN1(n1561), .IN2(n12), .QN(n1384) );
  NOR2X0 U937 ( .IN1(n1562), .IN2(n12), .QN(n1385) );
  NOR2X0 U938 ( .IN1(n1563), .IN2(n12), .QN(n1386) );
  NOR2X0 U939 ( .IN1(n1564), .IN2(n12), .QN(n1387) );
  NOR2X0 U940 ( .IN1(n1565), .IN2(n12), .QN(n1388) );
  NOR2X0 U941 ( .IN1(n1566), .IN2(n12), .QN(n1389) );
  NOR2X0 U942 ( .IN1(n80), .IN2(n1599), .QN(n1390) );
  NOR2X0 U943 ( .IN1(n78), .IN2(n12), .QN(n1391) );
  NOR2X0 U944 ( .IN1(n76), .IN2(n1599), .QN(n1392) );
  NOR2X0 U945 ( .IN1(n74), .IN2(n12), .QN(n1393) );
  NOR2X0 U946 ( .IN1(n1568), .IN2(n1599), .QN(n1394) );
  NOR2X0 U947 ( .IN1(n69), .IN2(n12), .QN(n1395) );
  NOR2X0 U948 ( .IN1(n67), .IN2(n1599), .QN(n1396) );
  NOR2X0 U949 ( .IN1(n65), .IN2(n1599), .QN(n1397) );
  NOR2X0 U950 ( .IN1(n1572), .IN2(n1599), .QN(n1398) );
  NOR2X0 U951 ( .IN1(n1573), .IN2(n1599), .QN(n1399) );
  NOR2X0 U952 ( .IN1(n59), .IN2(n1599), .QN(n1400) );
  NOR2X0 U953 ( .IN1(n57), .IN2(n1599), .QN(n1401) );
  NOR2X0 U954 ( .IN1(n55), .IN2(n1599), .QN(n1402) );
  NOR2X0 U955 ( .IN1(n53), .IN2(n1599), .QN(n1403) );
  NOR2X0 U956 ( .IN1(n51), .IN2(n1599), .QN(n1404) );
  NOR2X0 U957 ( .IN1(n1579), .IN2(n1599), .QN(n1405) );
  NOR2X0 U958 ( .IN1(n1555), .IN2(n1600), .QN(n1406) );
  NOR2X0 U959 ( .IN1(n1556), .IN2(n1600), .QN(n1407) );
  NOR2X0 U960 ( .IN1(n1557), .IN2(n1600), .QN(n1408) );
  NOR2X0 U961 ( .IN1(n1558), .IN2(n1600), .QN(n1409) );
  NOR2X0 U962 ( .IN1(n1559), .IN2(n1600), .QN(n1410) );
  NOR2X0 U963 ( .IN1(n1560), .IN2(n1600), .QN(n1411) );
  NOR2X0 U964 ( .IN1(n1561), .IN2(n1600), .QN(n1412) );
  NOR2X0 U965 ( .IN1(n1562), .IN2(n1600), .QN(n1413) );
  NOR2X0 U966 ( .IN1(n1563), .IN2(n1600), .QN(n1414) );
  NOR2X0 U967 ( .IN1(n1564), .IN2(n1600), .QN(n1415) );
  NOR2X0 U968 ( .IN1(n1565), .IN2(n1600), .QN(n1416) );
  NOR2X0 U969 ( .IN1(n1566), .IN2(n1600), .QN(n1417) );
  NOR2X0 U970 ( .IN1(n80), .IN2(n9), .QN(n1418) );
  NOR2X0 U971 ( .IN1(n78), .IN2(n9), .QN(n1419) );
  NOR2X0 U972 ( .IN1(n76), .IN2(n9), .QN(n1420) );
  NOR2X0 U973 ( .IN1(n1567), .IN2(n9), .QN(n1421) );
  NOR2X0 U974 ( .IN1(n1568), .IN2(n9), .QN(n1422) );
  NOR2X0 U975 ( .IN1(n69), .IN2(n9), .QN(n1423) );
  NOR2X0 U976 ( .IN1(n67), .IN2(n9), .QN(n1424) );
  NOR2X0 U977 ( .IN1(n65), .IN2(n9), .QN(n1425) );
  NOR2X0 U978 ( .IN1(n1572), .IN2(n9), .QN(n1426) );
  NOR2X0 U979 ( .IN1(n1573), .IN2(n9), .QN(n1427) );
  NOR2X0 U980 ( .IN1(n59), .IN2(n9), .QN(n1428) );
  NOR2X0 U981 ( .IN1(n57), .IN2(n9), .QN(n1429) );
  NOR2X0 U982 ( .IN1(n55), .IN2(n9), .QN(n1430) );
  NOR2X0 U983 ( .IN1(n53), .IN2(n9), .QN(n1431) );
  NOR2X0 U984 ( .IN1(n51), .IN2(n9), .QN(n1432) );
  NOR2X0 U985 ( .IN1(n1579), .IN2(n9), .QN(n1433) );
  NOR2X0 U986 ( .IN1(n93), .IN2(n8), .QN(n1434) );
  NOR2X0 U987 ( .IN1(n1555), .IN2(n8), .QN(n1435) );
  NOR2X0 U988 ( .IN1(n1556), .IN2(n8), .QN(n1436) );
  NOR2X0 U989 ( .IN1(n1557), .IN2(n8), .QN(n1437) );
  NOR2X0 U990 ( .IN1(n1558), .IN2(n8), .QN(n1438) );
  NOR2X0 U991 ( .IN1(n1559), .IN2(n8), .QN(n1439) );
  NOR2X0 U992 ( .IN1(n1560), .IN2(n8), .QN(n1440) );
  NOR2X0 U993 ( .IN1(n1561), .IN2(n8), .QN(n1441) );
  NOR2X0 U994 ( .IN1(n1562), .IN2(n8), .QN(n1442) );
  NOR2X0 U995 ( .IN1(n1563), .IN2(n8), .QN(n1443) );
  NOR2X0 U996 ( .IN1(n1564), .IN2(n8), .QN(n1444) );
  NOR2X0 U997 ( .IN1(n1565), .IN2(n8), .QN(n1445) );
  NOR2X0 U998 ( .IN1(n1566), .IN2(n8), .QN(n1446) );
  NOR2X0 U999 ( .IN1(n80), .IN2(n1601), .QN(n1447) );
  NOR2X0 U1000 ( .IN1(n78), .IN2(n8), .QN(n1448) );
  NOR2X0 U1001 ( .IN1(n76), .IN2(n1601), .QN(n1449) );
  NOR2X0 U1002 ( .IN1(n74), .IN2(n8), .QN(n1450) );
  NOR2X0 U1003 ( .IN1(n1568), .IN2(n1601), .QN(n1451) );
  NOR2X0 U1004 ( .IN1(n69), .IN2(n1601), .QN(n1452) );
  NOR2X0 U1005 ( .IN1(n67), .IN2(n1601), .QN(n1453) );
  NOR2X0 U1006 ( .IN1(n65), .IN2(n1601), .QN(n1454) );
  NOR2X0 U1007 ( .IN1(n1572), .IN2(n1601), .QN(n1455) );
  NOR2X0 U1008 ( .IN1(n1573), .IN2(n1601), .QN(n1456) );
  NOR2X0 U1009 ( .IN1(n59), .IN2(n1601), .QN(n1457) );
  NOR2X0 U1010 ( .IN1(n57), .IN2(n1601), .QN(n1458) );
  NOR2X0 U1011 ( .IN1(n55), .IN2(n1601), .QN(n1459) );
  NOR2X0 U1012 ( .IN1(n53), .IN2(n1601), .QN(n1460) );
  NOR2X0 U1013 ( .IN1(n51), .IN2(n1601), .QN(n1461) );
  NOR2X0 U1014 ( .IN1(n1579), .IN2(n1601), .QN(n1462) );
  NOR2X0 U1015 ( .IN1(n94), .IN2(n1602), .QN(n1463) );
  NOR2X0 U1016 ( .IN1(n93), .IN2(n1602), .QN(n1464) );
  NOR2X0 U1017 ( .IN1(n1555), .IN2(n1602), .QN(n1465) );
  NOR2X0 U1018 ( .IN1(n1556), .IN2(n1602), .QN(n1466) );
  NOR2X0 U1019 ( .IN1(n1557), .IN2(n1602), .QN(n1467) );
  NOR2X0 U1020 ( .IN1(n1558), .IN2(n1602), .QN(n1468) );
  NOR2X0 U1021 ( .IN1(n1559), .IN2(n1602), .QN(n1469) );
  NOR2X0 U1022 ( .IN1(n1560), .IN2(n1602), .QN(n1470) );
  NOR2X0 U1023 ( .IN1(n1561), .IN2(n1602), .QN(n1471) );
  NOR2X0 U1024 ( .IN1(n1562), .IN2(n1602), .QN(n1472) );
  NOR2X0 U1025 ( .IN1(n1563), .IN2(n1602), .QN(n1473) );
  NOR2X0 U1026 ( .IN1(n1564), .IN2(n1602), .QN(n1474) );
  NOR2X0 U1027 ( .IN1(n1565), .IN2(n1602), .QN(n1475) );
  NOR2X0 U1028 ( .IN1(n1566), .IN2(n1602), .QN(n1476) );
  NOR2X0 U1029 ( .IN1(n80), .IN2(n5), .QN(n1477) );
  NOR2X0 U1030 ( .IN1(n78), .IN2(n5), .QN(n1478) );
  NOR2X0 U1031 ( .IN1(n76), .IN2(n5), .QN(n1479) );
  NOR2X0 U1032 ( .IN1(n1567), .IN2(n5), .QN(n1480) );
  NOR2X0 U1033 ( .IN1(n1568), .IN2(n5), .QN(n1481) );
  NOR2X0 U1034 ( .IN1(n69), .IN2(n5), .QN(n1482) );
  NOR2X0 U1035 ( .IN1(n67), .IN2(n5), .QN(n1483) );
  NOR2X0 U1036 ( .IN1(n65), .IN2(n5), .QN(n1484) );
  NOR2X0 U1037 ( .IN1(n1572), .IN2(n5), .QN(n1485) );
  NOR2X0 U1038 ( .IN1(n1573), .IN2(n5), .QN(n1486) );
  NOR2X0 U1039 ( .IN1(n59), .IN2(n5), .QN(n1487) );
  NOR2X0 U1040 ( .IN1(n57), .IN2(n5), .QN(n1488) );
  NOR2X0 U1041 ( .IN1(n55), .IN2(n5), .QN(n1489) );
  NOR2X0 U1042 ( .IN1(n53), .IN2(n5), .QN(n1490) );
  NOR2X0 U1043 ( .IN1(n51), .IN2(n5), .QN(n1491) );
  NOR2X0 U1044 ( .IN1(n1579), .IN2(n5), .QN(n1492) );
  NOR2X0 U1045 ( .IN1(n95), .IN2(n1603), .QN(n1493) );
  NOR2X0 U1046 ( .IN1(n94), .IN2(n1603), .QN(n1494) );
  NOR2X0 U1047 ( .IN1(n93), .IN2(n1603), .QN(n1495) );
  NOR2X0 U1048 ( .IN1(n1555), .IN2(n1603), .QN(n1496) );
  NOR2X0 U1049 ( .IN1(n1556), .IN2(n1603), .QN(n1497) );
  NOR2X0 U1050 ( .IN1(n1557), .IN2(n1603), .QN(n1498) );
  NOR2X0 U1051 ( .IN1(n1558), .IN2(n1603), .QN(n1499) );
  NOR2X0 U1052 ( .IN1(n1559), .IN2(n1603), .QN(n1500) );
  NOR2X0 U1053 ( .IN1(n1560), .IN2(n1603), .QN(n1501) );
  NOR2X0 U1054 ( .IN1(n1561), .IN2(n1603), .QN(n1502) );
  NOR2X0 U1055 ( .IN1(n1562), .IN2(n1603), .QN(n1503) );
  NOR2X0 U1056 ( .IN1(n1563), .IN2(n1603), .QN(n1504) );
  NOR2X0 U1057 ( .IN1(n1564), .IN2(n1603), .QN(n1505) );
  NOR2X0 U1058 ( .IN1(n1565), .IN2(n1603), .QN(n1506) );
  NOR2X0 U1059 ( .IN1(n1566), .IN2(n1603), .QN(n1507) );
  NOR2X0 U1060 ( .IN1(n80), .IN2(n3), .QN(n1508) );
  NOR2X0 U1061 ( .IN1(n78), .IN2(n3), .QN(n1509) );
  NOR2X0 U1062 ( .IN1(n76), .IN2(n3), .QN(n1510) );
  NOR2X0 U1063 ( .IN1(n74), .IN2(n3), .QN(n1511) );
  NOR2X0 U1064 ( .IN1(n1568), .IN2(n3), .QN(n1512) );
  NOR2X0 U1065 ( .IN1(n69), .IN2(n3), .QN(n1513) );
  NOR2X0 U1066 ( .IN1(n67), .IN2(n3), .QN(n1514) );
  NOR2X0 U1067 ( .IN1(n65), .IN2(n3), .QN(n1515) );
  NOR2X0 U1068 ( .IN1(n1572), .IN2(n3), .QN(n1516) );
  NOR2X0 U1069 ( .IN1(n1573), .IN2(n3), .QN(n1517) );
  NOR2X0 U1070 ( .IN1(n59), .IN2(n3), .QN(n1518) );
  NOR2X0 U1071 ( .IN1(n57), .IN2(n3), .QN(n1519) );
  NOR2X0 U1072 ( .IN1(n55), .IN2(n3), .QN(n1520) );
  NOR2X0 U1073 ( .IN1(n53), .IN2(n3), .QN(n1521) );
  NOR2X0 U1074 ( .IN1(n51), .IN2(n3), .QN(n1522) );
  NOR2X0 U1075 ( .IN1(n1579), .IN2(n3), .QN(n1523) );
  NOR2X0 U1076 ( .IN1(n96), .IN2(n2), .QN(n1524) );
  NOR2X0 U1077 ( .IN1(n95), .IN2(n2), .QN(n1525) );
  NOR2X0 U1078 ( .IN1(n94), .IN2(n2), .QN(n1526) );
  NOR2X0 U1079 ( .IN1(n93), .IN2(n2), .QN(n1527) );
  NOR2X0 U1080 ( .IN1(n1555), .IN2(n2), .QN(n1528) );
  NOR2X0 U1081 ( .IN1(n1556), .IN2(n2), .QN(n1529) );
  NOR2X0 U1082 ( .IN1(n1557), .IN2(n2), .QN(n1530) );
  NOR2X0 U1083 ( .IN1(n1558), .IN2(n2), .QN(n1531) );
  NOR2X0 U1084 ( .IN1(n1559), .IN2(n2), .QN(n1532) );
  NOR2X0 U1085 ( .IN1(n1560), .IN2(n2), .QN(n1533) );
  NOR2X0 U1086 ( .IN1(n1561), .IN2(n2), .QN(n1534) );
  NOR2X0 U1087 ( .IN1(n1562), .IN2(n2), .QN(n1535) );
  NOR2X0 U1088 ( .IN1(n1563), .IN2(n2), .QN(n1536) );
  NOR2X0 U1089 ( .IN1(n1564), .IN2(n2), .QN(n1537) );
  NOR2X0 U1090 ( .IN1(n1565), .IN2(n2), .QN(n1538) );
  NOR2X0 U1091 ( .IN1(n1566), .IN2(n2), .QN(n1539) );
  NOR2X0 U1092 ( .IN1(n80), .IN2(n2), .QN(n1540) );
  NOR2X0 U1093 ( .IN1(n78), .IN2(n1604), .QN(n1541) );
  NOR2X0 U1094 ( .IN1(n76), .IN2(n1604), .QN(n1542) );
  NOR2X0 U1095 ( .IN1(n1567), .IN2(n1604), .QN(n1543) );
  NOR2X0 U1096 ( .IN1(n1568), .IN2(n1604), .QN(n1544) );
  NOR2X0 U1097 ( .IN1(n69), .IN2(n1604), .QN(n1545) );
  NOR2X0 U1098 ( .IN1(n67), .IN2(n1604), .QN(n1546) );
  NOR2X0 U1099 ( .IN1(n65), .IN2(n1604), .QN(n1547) );
  NOR2X0 U1100 ( .IN1(n1572), .IN2(n1604), .QN(n1548) );
  NOR2X0 U1101 ( .IN1(n1573), .IN2(n1604), .QN(n1549) );
  NOR2X0 U1102 ( .IN1(n59), .IN2(n1604), .QN(n1550) );
  NOR2X0 U1103 ( .IN1(n57), .IN2(n1604), .QN(n1551) );
  NOR2X0 U1104 ( .IN1(n55), .IN2(n1604), .QN(n1552) );
  NOR2X0 U1105 ( .IN1(n53), .IN2(n1604), .QN(n1553) );
  NOR2X0 U1106 ( .IN1(n51), .IN2(n1604), .QN(n1554) );
  NOR2X0 U1107 ( .IN1(n1579), .IN2(n1604), .QN(product[0]) );
  NBUFFX2 U1174 ( .INP(n1579), .Z(n50) );
  NBUFFX2 U1175 ( .INP(n1578), .Z(n51) );
  NBUFFX2 U1176 ( .INP(n1577), .Z(n53) );
  NBUFFX2 U1177 ( .INP(n1576), .Z(n55) );
  NBUFFX2 U1178 ( .INP(n1575), .Z(n57) );
  NBUFFX2 U1179 ( .INP(n1574), .Z(n59) );
  NBUFFX2 U1180 ( .INP(n1570), .Z(n67) );
  NBUFFX2 U1181 ( .INP(n1571), .Z(n65) );
  NBUFFX2 U1182 ( .INP(n1569), .Z(n69) );
  NBUFFX2 U1183 ( .INP(n1603), .Z(n3) );
  NBUFFX2 U1184 ( .INP(n1602), .Z(n5) );
  NBUFFX2 U1185 ( .INP(n1600), .Z(n9) );
  NBUFFX2 U1186 ( .INP(n1598), .Z(n13) );
  NBUFFX2 U1187 ( .INP(n1595), .Z(n19) );
  NBUFFX2 U1188 ( .INP(n1596), .Z(n17) );
  NBUFFX2 U1189 ( .INP(n1597), .Z(n15) );
  NBUFFX2 U1190 ( .INP(n1594), .Z(n21) );
  NBUFFX2 U1191 ( .INP(n1604), .Z(n2) );
  NBUFFX2 U1192 ( .INP(n1601), .Z(n8) );
  NBUFFX2 U1193 ( .INP(n1599), .Z(n12) );
  NBUFFX2 U1194 ( .INP(n1573), .Z(n62) );
  NBUFFX2 U1195 ( .INP(n1572), .Z(n64) );
  NBUFFX2 U1196 ( .INP(n1593), .Z(n24) );
  NBUFFX2 U1197 ( .INP(n1567), .Z(n74) );
  INVX0 U1198 ( .INP(b[0]), .ZN(n1579) );
  INVX0 U1199 ( .INP(b[1]), .ZN(n1578) );
  INVX0 U1200 ( .INP(b[2]), .ZN(n1577) );
  INVX0 U1201 ( .INP(b[3]), .ZN(n1576) );
  INVX0 U1202 ( .INP(b[4]), .ZN(n1575) );
  INVX0 U1203 ( .INP(b[16]), .ZN(n1566) );
  INVX0 U1204 ( .INP(a[16]), .ZN(n1591) );
  INVX0 U1205 ( .INP(b[17]), .ZN(n1565) );
  INVX0 U1206 ( .INP(a[17]), .ZN(n1590) );
  INVX0 U1207 ( .INP(b[18]), .ZN(n1564) );
  INVX0 U1208 ( .INP(a[18]), .ZN(n1589) );
  INVX0 U1209 ( .INP(b[19]), .ZN(n1563) );
  INVX0 U1210 ( .INP(a[19]), .ZN(n1588) );
  INVX0 U1211 ( .INP(b[20]), .ZN(n1562) );
  INVX0 U1212 ( .INP(a[20]), .ZN(n1587) );
  INVX0 U1213 ( .INP(b[21]), .ZN(n1561) );
  INVX0 U1214 ( .INP(a[21]), .ZN(n1586) );
  INVX0 U1215 ( .INP(b[22]), .ZN(n1560) );
  INVX0 U1216 ( .INP(a[22]), .ZN(n1585) );
  INVX0 U1217 ( .INP(b[23]), .ZN(n1559) );
  INVX0 U1218 ( .INP(a[23]), .ZN(n1584) );
  INVX0 U1219 ( .INP(b[24]), .ZN(n1558) );
  INVX0 U1220 ( .INP(a[24]), .ZN(n1583) );
  INVX0 U1221 ( .INP(b[25]), .ZN(n1557) );
  INVX0 U1222 ( .INP(a[25]), .ZN(n1582) );
  INVX0 U1223 ( .INP(b[26]), .ZN(n1556) );
  INVX0 U1224 ( .INP(a[26]), .ZN(n1581) );
  INVX0 U1225 ( .INP(b[27]), .ZN(n1555) );
  INVX0 U1226 ( .INP(a[27]), .ZN(n1580) );
  INVX0 U1227 ( .INP(b[5]), .ZN(n1574) );
  INVX0 U1228 ( .INP(b[7]), .ZN(n1572) );
  INVX0 U1229 ( .INP(b[6]), .ZN(n1573) );
  INVX0 U1230 ( .INP(b[9]), .ZN(n1570) );
  INVX0 U1231 ( .INP(b[8]), .ZN(n1571) );
  INVX0 U1232 ( .INP(b[10]), .ZN(n1569) );
  INVX0 U1233 ( .INP(b[11]), .ZN(n1568) );
  INVX0 U1234 ( .INP(b[12]), .ZN(n1567) );
  INVX0 U1235 ( .INP(a[1]), .ZN(n1603) );
  INVX0 U1236 ( .INP(a[2]), .ZN(n1602) );
  INVX0 U1237 ( .INP(a[3]), .ZN(n1601) );
  INVX0 U1238 ( .INP(a[4]), .ZN(n1600) );
  INVX0 U1239 ( .INP(a[5]), .ZN(n1599) );
  INVX0 U1240 ( .INP(a[6]), .ZN(n1598) );
  INVX0 U1241 ( .INP(a[9]), .ZN(n1595) );
  INVX0 U1242 ( .INP(a[8]), .ZN(n1596) );
  INVX0 U1243 ( .INP(a[7]), .ZN(n1597) );
  INVX0 U1244 ( .INP(a[10]), .ZN(n1594) );
  INVX0 U1245 ( .INP(a[11]), .ZN(n1593) );
  INVX0 U1246 ( .INP(a[12]), .ZN(n1592) );
  INVX0 U1247 ( .INP(b[13]), .ZN(n76) );
  INVX0 U1248 ( .INP(a[0]), .ZN(n1604) );
  INVX0 U1249 ( .INP(b[14]), .ZN(n78) );
  INVX0 U1250 ( .INP(b[15]), .ZN(n80) );
  INVX0 U1251 ( .INP(a[13]), .ZN(n28) );
  INVX0 U1252 ( .INP(a[14]), .ZN(n30) );
  INVX0 U1253 ( .INP(b[28]), .ZN(n93) );
  INVX0 U1254 ( .INP(a[31]), .ZN(n48) );
  INVX0 U1255 ( .INP(a[15]), .ZN(n32) );
  INVX0 U1256 ( .INP(b[29]), .ZN(n94) );
  INVX0 U1257 ( .INP(b[30]), .ZN(n95) );
  INVX0 U1258 ( .INP(b[31]), .ZN(n96) );
  INVX0 U1259 ( .INP(a[28]), .ZN(n45) );
  INVX0 U1260 ( .INP(a[29]), .ZN(n46) );
  INVX0 U1261 ( .INP(a[30]), .ZN(n47) );
endmodule


module thumb_DW_leftsh_3 ( A, SH, B );
  input [32:0] A;
  input [4:0] SH;
  output [32:0] B;
  wire   n1, n17, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163;

  MUX21X1 U1 ( .IN1(n57), .IN2(n41), .S(SH[4]), .Q(B[32]) );
  MUX21X1 U2 ( .IN1(n56), .IN2(n40), .S(SH[4]), .Q(B[31]) );
  MUX21X1 U3 ( .IN1(n55), .IN2(n39), .S(SH[4]), .Q(B[30]) );
  MUX21X1 U4 ( .IN1(n54), .IN2(n38), .S(SH[4]), .Q(B[29]) );
  MUX21X1 U5 ( .IN1(n53), .IN2(n37), .S(SH[4]), .Q(B[28]) );
  MUX21X1 U6 ( .IN1(n52), .IN2(n36), .S(SH[4]), .Q(B[27]) );
  MUX21X1 U7 ( .IN1(n51), .IN2(n35), .S(SH[4]), .Q(B[26]) );
  MUX21X1 U8 ( .IN1(n50), .IN2(n34), .S(SH[4]), .Q(B[25]) );
  MUX21X1 U9 ( .IN1(n49), .IN2(n33), .S(SH[4]), .Q(B[24]) );
  MUX21X1 U10 ( .IN1(n48), .IN2(n32), .S(SH[4]), .Q(B[23]) );
  MUX21X1 U11 ( .IN1(n47), .IN2(n31), .S(SH[4]), .Q(B[22]) );
  MUX21X1 U12 ( .IN1(n46), .IN2(n30), .S(SH[4]), .Q(B[21]) );
  MUX21X1 U13 ( .IN1(n45), .IN2(n29), .S(SH[4]), .Q(B[20]) );
  MUX21X1 U14 ( .IN1(n44), .IN2(n28), .S(SH[4]), .Q(B[19]) );
  MUX21X1 U15 ( .IN1(n43), .IN2(n27), .S(SH[4]), .Q(B[18]) );
  MUX21X1 U16 ( .IN1(n42), .IN2(n26), .S(SH[4]), .Q(B[17]) );
  MUX21X1 U17 ( .IN1(n41), .IN2(n25), .S(SH[4]), .Q(B[16]) );
  MUX21X1 U50 ( .IN1(n94), .IN2(n86), .S(SH[3]), .Q(n57) );
  MUX21X1 U51 ( .IN1(n93), .IN2(n85), .S(SH[3]), .Q(n56) );
  MUX21X1 U52 ( .IN1(n92), .IN2(n84), .S(SH[3]), .Q(n55) );
  MUX21X1 U53 ( .IN1(n91), .IN2(n83), .S(SH[3]), .Q(n54) );
  MUX21X1 U54 ( .IN1(n90), .IN2(n82), .S(SH[3]), .Q(n53) );
  MUX21X1 U55 ( .IN1(n89), .IN2(n81), .S(SH[3]), .Q(n52) );
  MUX21X1 U56 ( .IN1(n88), .IN2(n80), .S(SH[3]), .Q(n51) );
  MUX21X1 U57 ( .IN1(n87), .IN2(n79), .S(SH[3]), .Q(n50) );
  MUX21X1 U58 ( .IN1(n86), .IN2(n78), .S(SH[3]), .Q(n49) );
  MUX21X1 U59 ( .IN1(n85), .IN2(n77), .S(SH[3]), .Q(n48) );
  MUX21X1 U60 ( .IN1(n84), .IN2(n76), .S(SH[3]), .Q(n47) );
  MUX21X1 U61 ( .IN1(n83), .IN2(n75), .S(SH[3]), .Q(n46) );
  MUX21X1 U62 ( .IN1(n82), .IN2(n74), .S(SH[3]), .Q(n45) );
  MUX21X1 U63 ( .IN1(n81), .IN2(n73), .S(SH[3]), .Q(n44) );
  MUX21X1 U64 ( .IN1(n80), .IN2(n72), .S(SH[3]), .Q(n43) );
  MUX21X1 U65 ( .IN1(n79), .IN2(n71), .S(SH[3]), .Q(n42) );
  MUX21X1 U66 ( .IN1(n78), .IN2(n70), .S(SH[3]), .Q(n41) );
  MUX21X1 U67 ( .IN1(n77), .IN2(n69), .S(SH[3]), .Q(n40) );
  MUX21X1 U68 ( .IN1(n76), .IN2(n68), .S(SH[3]), .Q(n39) );
  MUX21X1 U69 ( .IN1(n75), .IN2(n67), .S(SH[3]), .Q(n38) );
  MUX21X1 U70 ( .IN1(n74), .IN2(n66), .S(SH[3]), .Q(n37) );
  MUX21X1 U71 ( .IN1(n73), .IN2(n65), .S(SH[3]), .Q(n36) );
  MUX21X1 U72 ( .IN1(n72), .IN2(n64), .S(SH[3]), .Q(n35) );
  MUX21X1 U73 ( .IN1(n71), .IN2(n63), .S(SH[3]), .Q(n34) );
  MUX21X1 U74 ( .IN1(n70), .IN2(n62), .S(SH[3]), .Q(n33) );
  MUX21X1 U91 ( .IN1(n129), .IN2(n125), .S(SH[2]), .Q(n94) );
  MUX21X1 U92 ( .IN1(n128), .IN2(n124), .S(SH[2]), .Q(n93) );
  MUX21X1 U93 ( .IN1(n127), .IN2(n123), .S(SH[2]), .Q(n92) );
  MUX21X1 U94 ( .IN1(n126), .IN2(n122), .S(SH[2]), .Q(n91) );
  MUX21X1 U95 ( .IN1(n125), .IN2(n121), .S(SH[2]), .Q(n90) );
  MUX21X1 U96 ( .IN1(n124), .IN2(n120), .S(SH[2]), .Q(n89) );
  MUX21X1 U97 ( .IN1(n123), .IN2(n119), .S(SH[2]), .Q(n88) );
  MUX21X1 U98 ( .IN1(n122), .IN2(n118), .S(SH[2]), .Q(n87) );
  MUX21X1 U99 ( .IN1(n121), .IN2(n117), .S(SH[2]), .Q(n86) );
  MUX21X1 U100 ( .IN1(n120), .IN2(n116), .S(SH[2]), .Q(n85) );
  MUX21X1 U101 ( .IN1(n119), .IN2(n115), .S(SH[2]), .Q(n84) );
  MUX21X1 U102 ( .IN1(n118), .IN2(n114), .S(SH[2]), .Q(n83) );
  MUX21X1 U103 ( .IN1(n117), .IN2(n113), .S(SH[2]), .Q(n82) );
  MUX21X1 U104 ( .IN1(n116), .IN2(n112), .S(SH[2]), .Q(n81) );
  MUX21X1 U105 ( .IN1(n115), .IN2(n111), .S(SH[2]), .Q(n80) );
  MUX21X1 U106 ( .IN1(n114), .IN2(n110), .S(SH[2]), .Q(n79) );
  MUX21X1 U107 ( .IN1(n113), .IN2(n109), .S(SH[2]), .Q(n78) );
  MUX21X1 U108 ( .IN1(n112), .IN2(n108), .S(SH[2]), .Q(n77) );
  MUX21X1 U109 ( .IN1(n111), .IN2(n107), .S(SH[2]), .Q(n76) );
  MUX21X1 U110 ( .IN1(n110), .IN2(n106), .S(SH[2]), .Q(n75) );
  MUX21X1 U111 ( .IN1(n109), .IN2(n105), .S(SH[2]), .Q(n74) );
  MUX21X1 U112 ( .IN1(n108), .IN2(n104), .S(SH[2]), .Q(n73) );
  MUX21X1 U113 ( .IN1(n107), .IN2(n103), .S(SH[2]), .Q(n72) );
  MUX21X1 U114 ( .IN1(n106), .IN2(n102), .S(SH[2]), .Q(n71) );
  MUX21X1 U115 ( .IN1(n105), .IN2(n101), .S(SH[2]), .Q(n70) );
  MUX21X1 U116 ( .IN1(n104), .IN2(n100), .S(SH[2]), .Q(n69) );
  MUX21X1 U117 ( .IN1(n103), .IN2(n99), .S(SH[2]), .Q(n68) );
  MUX21X1 U118 ( .IN1(n102), .IN2(n98), .S(SH[2]), .Q(n67) );
  MUX21X1 U119 ( .IN1(n101), .IN2(n97), .S(SH[2]), .Q(n66) );
  MUX21X1 U128 ( .IN1(n163), .IN2(n161), .S(SH[1]), .Q(n129) );
  MUX21X1 U129 ( .IN1(n162), .IN2(n160), .S(SH[1]), .Q(n128) );
  MUX21X1 U130 ( .IN1(n161), .IN2(n159), .S(SH[1]), .Q(n127) );
  MUX21X1 U131 ( .IN1(n160), .IN2(n158), .S(SH[1]), .Q(n126) );
  MUX21X1 U132 ( .IN1(n159), .IN2(n157), .S(SH[1]), .Q(n125) );
  MUX21X1 U133 ( .IN1(n158), .IN2(n156), .S(SH[1]), .Q(n124) );
  MUX21X1 U134 ( .IN1(n157), .IN2(n155), .S(SH[1]), .Q(n123) );
  MUX21X1 U135 ( .IN1(n156), .IN2(n154), .S(SH[1]), .Q(n122) );
  MUX21X1 U136 ( .IN1(n155), .IN2(n153), .S(SH[1]), .Q(n121) );
  MUX21X1 U137 ( .IN1(n154), .IN2(n152), .S(SH[1]), .Q(n120) );
  MUX21X1 U138 ( .IN1(n153), .IN2(n151), .S(SH[1]), .Q(n119) );
  MUX21X1 U139 ( .IN1(n152), .IN2(n150), .S(SH[1]), .Q(n118) );
  MUX21X1 U140 ( .IN1(n151), .IN2(n149), .S(SH[1]), .Q(n117) );
  MUX21X1 U141 ( .IN1(n150), .IN2(n148), .S(SH[1]), .Q(n116) );
  MUX21X1 U142 ( .IN1(n149), .IN2(n147), .S(SH[1]), .Q(n115) );
  MUX21X1 U143 ( .IN1(n148), .IN2(n146), .S(SH[1]), .Q(n114) );
  MUX21X1 U144 ( .IN1(n147), .IN2(n145), .S(SH[1]), .Q(n113) );
  MUX21X1 U145 ( .IN1(n146), .IN2(n144), .S(SH[1]), .Q(n112) );
  MUX21X1 U146 ( .IN1(n145), .IN2(n143), .S(SH[1]), .Q(n111) );
  MUX21X1 U147 ( .IN1(n144), .IN2(n142), .S(SH[1]), .Q(n110) );
  MUX21X1 U148 ( .IN1(n143), .IN2(n141), .S(SH[1]), .Q(n109) );
  MUX21X1 U149 ( .IN1(n142), .IN2(n140), .S(SH[1]), .Q(n108) );
  MUX21X1 U150 ( .IN1(n141), .IN2(n139), .S(SH[1]), .Q(n107) );
  MUX21X1 U151 ( .IN1(n140), .IN2(n138), .S(SH[1]), .Q(n106) );
  MUX21X1 U152 ( .IN1(n139), .IN2(n137), .S(SH[1]), .Q(n105) );
  MUX21X1 U153 ( .IN1(n138), .IN2(n136), .S(SH[1]), .Q(n104) );
  MUX21X1 U154 ( .IN1(n137), .IN2(n135), .S(SH[1]), .Q(n103) );
  MUX21X1 U155 ( .IN1(n136), .IN2(n134), .S(SH[1]), .Q(n102) );
  MUX21X1 U156 ( .IN1(n135), .IN2(n133), .S(SH[1]), .Q(n101) );
  MUX21X1 U157 ( .IN1(n134), .IN2(n132), .S(SH[1]), .Q(n100) );
  MUX21X1 U158 ( .IN1(n133), .IN2(n131), .S(SH[1]), .Q(n99) );
  AND2X1 U163 ( .IN1(SH[0]), .IN2(A[31]), .Q(n163) );
  MUX21X1 U164 ( .IN1(A[31]), .IN2(A[30]), .S(SH[0]), .Q(n162) );
  MUX21X1 U165 ( .IN1(A[30]), .IN2(A[29]), .S(SH[0]), .Q(n161) );
  MUX21X1 U166 ( .IN1(A[29]), .IN2(A[28]), .S(SH[0]), .Q(n160) );
  MUX21X1 U167 ( .IN1(A[28]), .IN2(A[27]), .S(SH[0]), .Q(n159) );
  MUX21X1 U168 ( .IN1(A[27]), .IN2(A[26]), .S(SH[0]), .Q(n158) );
  MUX21X1 U169 ( .IN1(A[26]), .IN2(A[25]), .S(SH[0]), .Q(n157) );
  MUX21X1 U170 ( .IN1(A[25]), .IN2(A[24]), .S(SH[0]), .Q(n156) );
  MUX21X1 U171 ( .IN1(A[24]), .IN2(A[23]), .S(SH[0]), .Q(n155) );
  MUX21X1 U172 ( .IN1(A[23]), .IN2(A[22]), .S(SH[0]), .Q(n154) );
  MUX21X1 U173 ( .IN1(A[22]), .IN2(A[21]), .S(SH[0]), .Q(n153) );
  MUX21X1 U174 ( .IN1(A[21]), .IN2(A[20]), .S(SH[0]), .Q(n152) );
  MUX21X1 U175 ( .IN1(A[20]), .IN2(A[19]), .S(SH[0]), .Q(n151) );
  MUX21X1 U176 ( .IN1(A[19]), .IN2(A[18]), .S(SH[0]), .Q(n150) );
  MUX21X1 U177 ( .IN1(A[18]), .IN2(A[17]), .S(SH[0]), .Q(n149) );
  MUX21X1 U178 ( .IN1(A[17]), .IN2(A[16]), .S(SH[0]), .Q(n148) );
  MUX21X1 U179 ( .IN1(A[16]), .IN2(A[15]), .S(SH[0]), .Q(n147) );
  MUX21X1 U180 ( .IN1(A[15]), .IN2(A[14]), .S(SH[0]), .Q(n146) );
  MUX21X1 U181 ( .IN1(A[14]), .IN2(A[13]), .S(SH[0]), .Q(n145) );
  MUX21X1 U182 ( .IN1(A[13]), .IN2(A[12]), .S(SH[0]), .Q(n144) );
  MUX21X1 U183 ( .IN1(A[12]), .IN2(A[11]), .S(SH[0]), .Q(n143) );
  MUX21X1 U184 ( .IN1(A[11]), .IN2(A[10]), .S(SH[0]), .Q(n142) );
  MUX21X1 U185 ( .IN1(A[10]), .IN2(A[9]), .S(SH[0]), .Q(n141) );
  MUX21X1 U186 ( .IN1(A[9]), .IN2(A[8]), .S(SH[0]), .Q(n140) );
  MUX21X1 U187 ( .IN1(A[8]), .IN2(A[7]), .S(SH[0]), .Q(n139) );
  MUX21X1 U188 ( .IN1(A[7]), .IN2(A[6]), .S(SH[0]), .Q(n138) );
  MUX21X1 U189 ( .IN1(A[6]), .IN2(A[5]), .S(SH[0]), .Q(n137) );
  MUX21X1 U190 ( .IN1(A[5]), .IN2(A[4]), .S(SH[0]), .Q(n136) );
  MUX21X1 U191 ( .IN1(A[4]), .IN2(A[3]), .S(SH[0]), .Q(n135) );
  MUX21X1 U192 ( .IN1(A[3]), .IN2(A[2]), .S(SH[0]), .Q(n134) );
  MUX21X1 U193 ( .IN1(A[2]), .IN2(A[1]), .S(SH[0]), .Q(n133) );
  MUX21X1 U194 ( .IN1(A[1]), .IN2(A[0]), .S(SH[0]), .Q(n132) );
  AND2X1 U200 ( .IN1(A[0]), .IN2(n130), .Q(n131) );
  AND2X1 U201 ( .IN1(n33), .IN2(n1), .Q(B[8]) );
  AND2X1 U202 ( .IN1(n26), .IN2(n1), .Q(B[1]) );
  AND2X1 U203 ( .IN1(n40), .IN2(n1), .Q(B[15]) );
  AND2X1 U204 ( .IN1(n39), .IN2(n1), .Q(B[14]) );
  AND2X1 U205 ( .IN1(n38), .IN2(n1), .Q(B[13]) );
  AND2X1 U206 ( .IN1(n36), .IN2(n1), .Q(B[11]) );
  AND2X1 U207 ( .IN1(n35), .IN2(n1), .Q(B[10]) );
  AND2X1 U208 ( .IN1(n34), .IN2(n1), .Q(B[9]) );
  AND2X1 U209 ( .IN1(n32), .IN2(n1), .Q(B[7]) );
  AND2X1 U210 ( .IN1(n31), .IN2(n1), .Q(B[6]) );
  AND2X1 U211 ( .IN1(n30), .IN2(n1), .Q(B[5]) );
  AND2X1 U212 ( .IN1(n29), .IN2(n1), .Q(B[4]) );
  AND2X1 U213 ( .IN1(n28), .IN2(n1), .Q(B[3]) );
  AND2X1 U214 ( .IN1(n27), .IN2(n1), .Q(B[2]) );
  AND2X1 U215 ( .IN1(n25), .IN2(n1), .Q(B[0]) );
  AND2X1 U216 ( .IN1(n37), .IN2(n1), .Q(B[12]) );
  AND2X1 U217 ( .IN1(n69), .IN2(n17), .Q(n32) );
  AND2X1 U218 ( .IN1(n68), .IN2(n17), .Q(n31) );
  AND2X1 U219 ( .IN1(n67), .IN2(n17), .Q(n30) );
  AND2X1 U220 ( .IN1(n66), .IN2(n17), .Q(n29) );
  AND2X1 U221 ( .IN1(n65), .IN2(n17), .Q(n28) );
  AND2X1 U222 ( .IN1(n64), .IN2(n17), .Q(n27) );
  AND2X1 U223 ( .IN1(n63), .IN2(n17), .Q(n26) );
  AND2X1 U224 ( .IN1(n62), .IN2(n17), .Q(n25) );
  AND2X1 U225 ( .IN1(n100), .IN2(n58), .Q(n65) );
  AND2X1 U226 ( .IN1(n99), .IN2(n58), .Q(n64) );
  AND2X1 U227 ( .IN1(n98), .IN2(n58), .Q(n63) );
  AND2X1 U228 ( .IN1(n97), .IN2(n58), .Q(n62) );
  AND2X1 U229 ( .IN1(n132), .IN2(n95), .Q(n98) );
  AND2X1 U230 ( .IN1(n131), .IN2(n95), .Q(n97) );
  INVX0 U231 ( .INP(SH[4]), .ZN(n1) );
  INVX0 U232 ( .INP(SH[3]), .ZN(n17) );
  INVX0 U233 ( .INP(SH[2]), .ZN(n58) );
  INVX0 U234 ( .INP(SH[1]), .ZN(n95) );
  INVX0 U235 ( .INP(SH[0]), .ZN(n130) );
endmodule


module thumb_DW_rightsh_4 ( A, DATA_TC, SH, B );
  input [32:0] A;
  input [4:0] SH;
  output [32:0] B;
  input DATA_TC;
  wire   n1, n17, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163;

  MUX21X1 U33 ( .IN1(n41), .IN2(n57), .S(SH[4]), .Q(B[16]) );
  MUX21X1 U34 ( .IN1(n40), .IN2(n56), .S(SH[4]), .Q(B[15]) );
  MUX21X1 U35 ( .IN1(n39), .IN2(n55), .S(SH[4]), .Q(B[14]) );
  MUX21X1 U36 ( .IN1(n38), .IN2(n54), .S(SH[4]), .Q(B[13]) );
  MUX21X1 U37 ( .IN1(n37), .IN2(n53), .S(SH[4]), .Q(B[12]) );
  MUX21X1 U38 ( .IN1(n36), .IN2(n52), .S(SH[4]), .Q(B[11]) );
  MUX21X1 U39 ( .IN1(n35), .IN2(n51), .S(SH[4]), .Q(B[10]) );
  MUX21X1 U40 ( .IN1(n34), .IN2(n50), .S(SH[4]), .Q(B[9]) );
  MUX21X1 U41 ( .IN1(n33), .IN2(n49), .S(SH[4]), .Q(B[8]) );
  MUX21X1 U42 ( .IN1(n32), .IN2(n48), .S(SH[4]), .Q(B[7]) );
  MUX21X1 U43 ( .IN1(n31), .IN2(n47), .S(SH[4]), .Q(B[6]) );
  MUX21X1 U44 ( .IN1(n30), .IN2(n46), .S(SH[4]), .Q(B[5]) );
  MUX21X1 U45 ( .IN1(n29), .IN2(n45), .S(SH[4]), .Q(B[4]) );
  MUX21X1 U46 ( .IN1(n28), .IN2(n44), .S(SH[4]), .Q(B[3]) );
  MUX21X1 U47 ( .IN1(n27), .IN2(n43), .S(SH[4]), .Q(B[2]) );
  MUX21X1 U48 ( .IN1(n26), .IN2(n42), .S(SH[4]), .Q(B[1]) );
  MUX21X1 U49 ( .IN1(n25), .IN2(n41), .S(SH[4]), .Q(B[0]) );
  MUX21X1 U66 ( .IN1(n86), .IN2(n94), .S(SH[3]), .Q(n49) );
  MUX21X1 U67 ( .IN1(n85), .IN2(n93), .S(SH[3]), .Q(n48) );
  MUX21X1 U68 ( .IN1(n84), .IN2(n92), .S(SH[3]), .Q(n47) );
  MUX21X1 U69 ( .IN1(n83), .IN2(n91), .S(SH[3]), .Q(n46) );
  MUX21X1 U70 ( .IN1(n82), .IN2(n90), .S(SH[3]), .Q(n45) );
  MUX21X1 U71 ( .IN1(n81), .IN2(n89), .S(SH[3]), .Q(n44) );
  MUX21X1 U72 ( .IN1(n80), .IN2(n88), .S(SH[3]), .Q(n43) );
  MUX21X1 U73 ( .IN1(n79), .IN2(n87), .S(SH[3]), .Q(n42) );
  MUX21X1 U74 ( .IN1(n78), .IN2(n86), .S(SH[3]), .Q(n41) );
  MUX21X1 U75 ( .IN1(n77), .IN2(n85), .S(SH[3]), .Q(n40) );
  MUX21X1 U76 ( .IN1(n76), .IN2(n84), .S(SH[3]), .Q(n39) );
  MUX21X1 U77 ( .IN1(n75), .IN2(n83), .S(SH[3]), .Q(n38) );
  MUX21X1 U78 ( .IN1(n74), .IN2(n82), .S(SH[3]), .Q(n37) );
  MUX21X1 U79 ( .IN1(n73), .IN2(n81), .S(SH[3]), .Q(n36) );
  MUX21X1 U80 ( .IN1(n72), .IN2(n80), .S(SH[3]), .Q(n35) );
  MUX21X1 U81 ( .IN1(n71), .IN2(n79), .S(SH[3]), .Q(n34) );
  MUX21X1 U82 ( .IN1(n70), .IN2(n78), .S(SH[3]), .Q(n33) );
  MUX21X1 U83 ( .IN1(n69), .IN2(n77), .S(SH[3]), .Q(n32) );
  MUX21X1 U84 ( .IN1(n68), .IN2(n76), .S(SH[3]), .Q(n31) );
  MUX21X1 U85 ( .IN1(n67), .IN2(n75), .S(SH[3]), .Q(n30) );
  MUX21X1 U86 ( .IN1(n66), .IN2(n74), .S(SH[3]), .Q(n29) );
  MUX21X1 U87 ( .IN1(n65), .IN2(n73), .S(SH[3]), .Q(n28) );
  MUX21X1 U88 ( .IN1(n64), .IN2(n72), .S(SH[3]), .Q(n27) );
  MUX21X1 U89 ( .IN1(n63), .IN2(n71), .S(SH[3]), .Q(n26) );
  MUX21X1 U90 ( .IN1(n62), .IN2(n70), .S(SH[3]), .Q(n25) );
  MUX21X1 U99 ( .IN1(n125), .IN2(n129), .S(SH[2]), .Q(n90) );
  MUX21X1 U100 ( .IN1(n124), .IN2(n128), .S(SH[2]), .Q(n89) );
  MUX21X1 U101 ( .IN1(n123), .IN2(n127), .S(SH[2]), .Q(n88) );
  MUX21X1 U102 ( .IN1(n122), .IN2(n126), .S(SH[2]), .Q(n87) );
  MUX21X1 U103 ( .IN1(n121), .IN2(n125), .S(SH[2]), .Q(n86) );
  MUX21X1 U104 ( .IN1(n120), .IN2(n124), .S(SH[2]), .Q(n85) );
  MUX21X1 U105 ( .IN1(n119), .IN2(n123), .S(SH[2]), .Q(n84) );
  MUX21X1 U106 ( .IN1(n118), .IN2(n122), .S(SH[2]), .Q(n83) );
  MUX21X1 U107 ( .IN1(n117), .IN2(n121), .S(SH[2]), .Q(n82) );
  MUX21X1 U108 ( .IN1(n116), .IN2(n120), .S(SH[2]), .Q(n81) );
  MUX21X1 U109 ( .IN1(n115), .IN2(n119), .S(SH[2]), .Q(n80) );
  MUX21X1 U110 ( .IN1(n114), .IN2(n118), .S(SH[2]), .Q(n79) );
  MUX21X1 U111 ( .IN1(n113), .IN2(n117), .S(SH[2]), .Q(n78) );
  MUX21X1 U112 ( .IN1(n112), .IN2(n116), .S(SH[2]), .Q(n77) );
  MUX21X1 U113 ( .IN1(n111), .IN2(n115), .S(SH[2]), .Q(n76) );
  MUX21X1 U114 ( .IN1(n110), .IN2(n114), .S(SH[2]), .Q(n75) );
  MUX21X1 U115 ( .IN1(n109), .IN2(n113), .S(SH[2]), .Q(n74) );
  MUX21X1 U116 ( .IN1(n108), .IN2(n112), .S(SH[2]), .Q(n73) );
  MUX21X1 U117 ( .IN1(n107), .IN2(n111), .S(SH[2]), .Q(n72) );
  MUX21X1 U118 ( .IN1(n106), .IN2(n110), .S(SH[2]), .Q(n71) );
  MUX21X1 U119 ( .IN1(n105), .IN2(n109), .S(SH[2]), .Q(n70) );
  MUX21X1 U120 ( .IN1(n104), .IN2(n108), .S(SH[2]), .Q(n69) );
  MUX21X1 U121 ( .IN1(n103), .IN2(n107), .S(SH[2]), .Q(n68) );
  MUX21X1 U122 ( .IN1(n102), .IN2(n106), .S(SH[2]), .Q(n67) );
  MUX21X1 U123 ( .IN1(n101), .IN2(n105), .S(SH[2]), .Q(n66) );
  MUX21X1 U124 ( .IN1(n100), .IN2(n104), .S(SH[2]), .Q(n65) );
  MUX21X1 U125 ( .IN1(n99), .IN2(n103), .S(SH[2]), .Q(n64) );
  MUX21X1 U126 ( .IN1(n98), .IN2(n102), .S(SH[2]), .Q(n63) );
  MUX21X1 U127 ( .IN1(n97), .IN2(n101), .S(SH[2]), .Q(n62) );
  MUX21X1 U132 ( .IN1(n161), .IN2(n163), .S(SH[1]), .Q(n127) );
  MUX21X1 U133 ( .IN1(n160), .IN2(n162), .S(SH[1]), .Q(n126) );
  MUX21X1 U134 ( .IN1(n159), .IN2(n161), .S(SH[1]), .Q(n125) );
  MUX21X1 U135 ( .IN1(n158), .IN2(n160), .S(SH[1]), .Q(n124) );
  MUX21X1 U136 ( .IN1(n157), .IN2(n159), .S(SH[1]), .Q(n123) );
  MUX21X1 U137 ( .IN1(n156), .IN2(n158), .S(SH[1]), .Q(n122) );
  MUX21X1 U138 ( .IN1(n155), .IN2(n157), .S(SH[1]), .Q(n121) );
  MUX21X1 U139 ( .IN1(n154), .IN2(n156), .S(SH[1]), .Q(n120) );
  MUX21X1 U140 ( .IN1(n153), .IN2(n155), .S(SH[1]), .Q(n119) );
  MUX21X1 U141 ( .IN1(n152), .IN2(n154), .S(SH[1]), .Q(n118) );
  MUX21X1 U142 ( .IN1(n151), .IN2(n153), .S(SH[1]), .Q(n117) );
  MUX21X1 U143 ( .IN1(n150), .IN2(n152), .S(SH[1]), .Q(n116) );
  MUX21X1 U144 ( .IN1(n149), .IN2(n151), .S(SH[1]), .Q(n115) );
  MUX21X1 U145 ( .IN1(n148), .IN2(n150), .S(SH[1]), .Q(n114) );
  MUX21X1 U146 ( .IN1(n147), .IN2(n149), .S(SH[1]), .Q(n113) );
  MUX21X1 U147 ( .IN1(n146), .IN2(n148), .S(SH[1]), .Q(n112) );
  MUX21X1 U148 ( .IN1(n145), .IN2(n147), .S(SH[1]), .Q(n111) );
  MUX21X1 U149 ( .IN1(n144), .IN2(n146), .S(SH[1]), .Q(n110) );
  MUX21X1 U150 ( .IN1(n143), .IN2(n145), .S(SH[1]), .Q(n109) );
  MUX21X1 U151 ( .IN1(n142), .IN2(n144), .S(SH[1]), .Q(n108) );
  MUX21X1 U152 ( .IN1(n141), .IN2(n143), .S(SH[1]), .Q(n107) );
  MUX21X1 U153 ( .IN1(n140), .IN2(n142), .S(SH[1]), .Q(n106) );
  MUX21X1 U154 ( .IN1(n139), .IN2(n141), .S(SH[1]), .Q(n105) );
  MUX21X1 U155 ( .IN1(n138), .IN2(n140), .S(SH[1]), .Q(n104) );
  MUX21X1 U156 ( .IN1(n137), .IN2(n139), .S(SH[1]), .Q(n103) );
  MUX21X1 U157 ( .IN1(n136), .IN2(n138), .S(SH[1]), .Q(n102) );
  MUX21X1 U158 ( .IN1(n135), .IN2(n137), .S(SH[1]), .Q(n101) );
  MUX21X1 U159 ( .IN1(n134), .IN2(n136), .S(SH[1]), .Q(n100) );
  MUX21X1 U160 ( .IN1(n133), .IN2(n135), .S(SH[1]), .Q(n99) );
  MUX21X1 U161 ( .IN1(n132), .IN2(n134), .S(SH[1]), .Q(n98) );
  MUX21X1 U162 ( .IN1(n131), .IN2(n133), .S(SH[1]), .Q(n97) );
  MUX21X1 U165 ( .IN1(A[31]), .IN2(A[32]), .S(SH[0]), .Q(n162) );
  MUX21X1 U166 ( .IN1(A[30]), .IN2(A[31]), .S(SH[0]), .Q(n161) );
  MUX21X1 U167 ( .IN1(A[29]), .IN2(A[30]), .S(SH[0]), .Q(n160) );
  MUX21X1 U168 ( .IN1(A[28]), .IN2(A[29]), .S(SH[0]), .Q(n159) );
  MUX21X1 U169 ( .IN1(A[27]), .IN2(A[28]), .S(SH[0]), .Q(n158) );
  MUX21X1 U170 ( .IN1(A[26]), .IN2(A[27]), .S(SH[0]), .Q(n157) );
  MUX21X1 U171 ( .IN1(A[25]), .IN2(A[26]), .S(SH[0]), .Q(n156) );
  MUX21X1 U172 ( .IN1(A[24]), .IN2(A[25]), .S(SH[0]), .Q(n155) );
  MUX21X1 U173 ( .IN1(A[23]), .IN2(A[24]), .S(SH[0]), .Q(n154) );
  MUX21X1 U174 ( .IN1(A[22]), .IN2(A[23]), .S(SH[0]), .Q(n153) );
  MUX21X1 U175 ( .IN1(A[21]), .IN2(A[22]), .S(SH[0]), .Q(n152) );
  MUX21X1 U176 ( .IN1(A[20]), .IN2(A[21]), .S(SH[0]), .Q(n151) );
  MUX21X1 U177 ( .IN1(A[19]), .IN2(A[20]), .S(SH[0]), .Q(n150) );
  MUX21X1 U178 ( .IN1(A[18]), .IN2(A[19]), .S(SH[0]), .Q(n149) );
  MUX21X1 U179 ( .IN1(A[17]), .IN2(A[18]), .S(SH[0]), .Q(n148) );
  MUX21X1 U180 ( .IN1(A[16]), .IN2(A[17]), .S(SH[0]), .Q(n147) );
  MUX21X1 U181 ( .IN1(A[15]), .IN2(A[16]), .S(SH[0]), .Q(n146) );
  MUX21X1 U182 ( .IN1(A[14]), .IN2(A[15]), .S(SH[0]), .Q(n145) );
  MUX21X1 U183 ( .IN1(A[13]), .IN2(A[14]), .S(SH[0]), .Q(n144) );
  MUX21X1 U184 ( .IN1(A[12]), .IN2(A[13]), .S(SH[0]), .Q(n143) );
  MUX21X1 U185 ( .IN1(A[11]), .IN2(A[12]), .S(SH[0]), .Q(n142) );
  MUX21X1 U186 ( .IN1(A[10]), .IN2(A[11]), .S(SH[0]), .Q(n141) );
  MUX21X1 U187 ( .IN1(A[9]), .IN2(A[10]), .S(SH[0]), .Q(n140) );
  MUX21X1 U188 ( .IN1(A[8]), .IN2(A[9]), .S(SH[0]), .Q(n139) );
  MUX21X1 U189 ( .IN1(A[7]), .IN2(A[8]), .S(SH[0]), .Q(n138) );
  MUX21X1 U190 ( .IN1(A[6]), .IN2(A[7]), .S(SH[0]), .Q(n137) );
  MUX21X1 U191 ( .IN1(A[5]), .IN2(A[6]), .S(SH[0]), .Q(n136) );
  MUX21X1 U192 ( .IN1(A[4]), .IN2(A[5]), .S(SH[0]), .Q(n135) );
  MUX21X1 U193 ( .IN1(A[3]), .IN2(A[4]), .S(SH[0]), .Q(n134) );
  MUX21X1 U194 ( .IN1(A[2]), .IN2(A[3]), .S(SH[0]), .Q(n133) );
  MUX21X1 U195 ( .IN1(A[1]), .IN2(A[2]), .S(SH[0]), .Q(n132) );
  AND2X1 U196 ( .IN1(SH[0]), .IN2(A[1]), .Q(n131) );
  AND2X1 U200 ( .IN1(n56), .IN2(n1), .Q(B[31]) );
  AND2X1 U201 ( .IN1(n55), .IN2(n1), .Q(B[30]) );
  AND2X1 U202 ( .IN1(n54), .IN2(n1), .Q(B[29]) );
  AND2X1 U203 ( .IN1(n53), .IN2(n1), .Q(B[28]) );
  AND2X1 U204 ( .IN1(n52), .IN2(n1), .Q(B[27]) );
  AND2X1 U205 ( .IN1(n51), .IN2(n1), .Q(B[26]) );
  AND2X1 U206 ( .IN1(n50), .IN2(n1), .Q(B[25]) );
  AND2X1 U207 ( .IN1(n49), .IN2(n1), .Q(B[24]) );
  AND2X1 U208 ( .IN1(n48), .IN2(n1), .Q(B[23]) );
  AND2X1 U209 ( .IN1(n47), .IN2(n1), .Q(B[22]) );
  AND2X1 U210 ( .IN1(n46), .IN2(n1), .Q(B[21]) );
  AND2X1 U211 ( .IN1(n44), .IN2(n1), .Q(B[19]) );
  AND2X1 U212 ( .IN1(n43), .IN2(n1), .Q(B[18]) );
  AND2X1 U213 ( .IN1(n42), .IN2(n1), .Q(B[17]) );
  AND2X1 U214 ( .IN1(n45), .IN2(n1), .Q(B[20]) );
  AND2X1 U215 ( .IN1(n94), .IN2(n17), .Q(n57) );
  AND2X1 U216 ( .IN1(n93), .IN2(n17), .Q(n56) );
  AND2X1 U217 ( .IN1(n92), .IN2(n17), .Q(n55) );
  AND2X1 U218 ( .IN1(n91), .IN2(n17), .Q(n54) );
  AND2X1 U219 ( .IN1(n90), .IN2(n17), .Q(n53) );
  AND2X1 U220 ( .IN1(n89), .IN2(n17), .Q(n52) );
  AND2X1 U221 ( .IN1(n88), .IN2(n17), .Q(n51) );
  AND2X1 U222 ( .IN1(n87), .IN2(n17), .Q(n50) );
  AND2X1 U223 ( .IN1(n129), .IN2(n58), .Q(n94) );
  AND2X1 U224 ( .IN1(n128), .IN2(n58), .Q(n93) );
  AND2X1 U225 ( .IN1(n127), .IN2(n58), .Q(n92) );
  AND2X1 U226 ( .IN1(n126), .IN2(n58), .Q(n91) );
  AND2X1 U227 ( .IN1(n163), .IN2(n95), .Q(n129) );
  AND2X1 U228 ( .IN1(n162), .IN2(n95), .Q(n128) );
  AND2X1 U229 ( .IN1(n57), .IN2(n1), .Q(B[32]) );
  INVX0 U230 ( .INP(SH[4]), .ZN(n1) );
  INVX0 U231 ( .INP(SH[3]), .ZN(n17) );
  INVX0 U232 ( .INP(SH[2]), .ZN(n58) );
  INVX0 U233 ( .INP(SH[1]), .ZN(n95) );
  AND2X1 U234 ( .IN1(A[32]), .IN2(n130), .Q(n163) );
  INVX0 U235 ( .INP(SH[0]), .ZN(n130) );
endmodule


module thumb_DW_rightsh_5 ( A, DATA_TC, SH, B );
  input [32:0] A;
  input [7:0] SH;
  output [32:0] B;
  input DATA_TC;
  wire   n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n44, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n81, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n118, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n155, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n191, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n307;

  AND2X1 U4 ( .IN1(n41), .IN2(n307), .Q(B[32]) );
  AND2X1 U5 ( .IN1(n40), .IN2(n307), .Q(B[31]) );
  AND2X1 U6 ( .IN1(n39), .IN2(n307), .Q(B[30]) );
  AND2X1 U7 ( .IN1(n38), .IN2(n307), .Q(B[29]) );
  AND2X1 U8 ( .IN1(n37), .IN2(n307), .Q(B[28]) );
  AND2X1 U9 ( .IN1(n36), .IN2(n307), .Q(B[27]) );
  AND2X1 U10 ( .IN1(n35), .IN2(n307), .Q(B[26]) );
  AND2X1 U11 ( .IN1(n34), .IN2(n307), .Q(B[25]) );
  AND2X1 U12 ( .IN1(n33), .IN2(n307), .Q(B[24]) );
  AND2X1 U13 ( .IN1(n32), .IN2(n307), .Q(B[23]) );
  AND2X1 U14 ( .IN1(n31), .IN2(n307), .Q(B[22]) );
  AND2X1 U15 ( .IN1(n30), .IN2(n307), .Q(B[21]) );
  AND2X1 U16 ( .IN1(n29), .IN2(n307), .Q(B[20]) );
  AND2X1 U17 ( .IN1(n28), .IN2(n307), .Q(B[19]) );
  AND2X1 U18 ( .IN1(n27), .IN2(n307), .Q(B[18]) );
  AND2X1 U19 ( .IN1(n26), .IN2(n307), .Q(B[17]) );
  AND2X1 U20 ( .IN1(n25), .IN2(n307), .Q(B[16]) );
  AND2X1 U21 ( .IN1(n24), .IN2(n307), .Q(B[15]) );
  AND2X1 U22 ( .IN1(n23), .IN2(n307), .Q(B[14]) );
  AND2X1 U23 ( .IN1(n22), .IN2(n307), .Q(B[13]) );
  AND2X1 U24 ( .IN1(n21), .IN2(n307), .Q(B[12]) );
  AND2X1 U25 ( .IN1(n20), .IN2(n307), .Q(B[11]) );
  AND2X1 U26 ( .IN1(n19), .IN2(n307), .Q(B[10]) );
  AND2X1 U27 ( .IN1(n18), .IN2(n307), .Q(B[9]) );
  AND2X1 U28 ( .IN1(n17), .IN2(n307), .Q(B[8]) );
  AND2X1 U29 ( .IN1(n16), .IN2(n307), .Q(B[7]) );
  AND2X1 U30 ( .IN1(n15), .IN2(n307), .Q(B[6]) );
  AND2X1 U31 ( .IN1(n14), .IN2(n307), .Q(B[5]) );
  AND2X1 U32 ( .IN1(n13), .IN2(n307), .Q(B[4]) );
  AND2X1 U33 ( .IN1(n12), .IN2(n307), .Q(B[3]) );
  AND2X1 U34 ( .IN1(n11), .IN2(n307), .Q(B[2]) );
  AND2X1 U35 ( .IN1(n10), .IN2(n307), .Q(B[1]) );
  AND2X1 U36 ( .IN1(n9), .IN2(n307), .Q(B[0]) );
  AND2X1 U41 ( .IN1(n78), .IN2(n7), .Q(n41) );
  AND2X1 U42 ( .IN1(n77), .IN2(n7), .Q(n40) );
  AND2X1 U43 ( .IN1(n76), .IN2(n7), .Q(n39) );
  AND2X1 U44 ( .IN1(n75), .IN2(n7), .Q(n38) );
  AND2X1 U45 ( .IN1(n74), .IN2(n7), .Q(n37) );
  AND2X1 U46 ( .IN1(n73), .IN2(n7), .Q(n36) );
  AND2X1 U47 ( .IN1(n72), .IN2(n7), .Q(n35) );
  AND2X1 U48 ( .IN1(n71), .IN2(n7), .Q(n34) );
  AND2X1 U49 ( .IN1(n70), .IN2(n7), .Q(n33) );
  AND2X1 U50 ( .IN1(n69), .IN2(n7), .Q(n32) );
  AND2X1 U51 ( .IN1(n68), .IN2(n7), .Q(n31) );
  AND2X1 U52 ( .IN1(n67), .IN2(n7), .Q(n30) );
  AND2X1 U53 ( .IN1(n66), .IN2(n7), .Q(n29) );
  AND2X1 U54 ( .IN1(n65), .IN2(n7), .Q(n28) );
  AND2X1 U55 ( .IN1(n64), .IN2(n7), .Q(n27) );
  AND2X1 U56 ( .IN1(n63), .IN2(n7), .Q(n26) );
  AND2X1 U57 ( .IN1(n62), .IN2(n7), .Q(n25) );
  AND2X1 U58 ( .IN1(n61), .IN2(n7), .Q(n24) );
  AND2X1 U59 ( .IN1(n60), .IN2(n7), .Q(n23) );
  AND2X1 U60 ( .IN1(n59), .IN2(n7), .Q(n22) );
  AND2X1 U61 ( .IN1(n58), .IN2(n7), .Q(n21) );
  AND2X1 U62 ( .IN1(n57), .IN2(n7), .Q(n20) );
  AND2X1 U63 ( .IN1(n56), .IN2(n7), .Q(n19) );
  AND2X1 U64 ( .IN1(n55), .IN2(n7), .Q(n18) );
  AND2X1 U65 ( .IN1(n54), .IN2(n7), .Q(n17) );
  AND2X1 U66 ( .IN1(n53), .IN2(n7), .Q(n16) );
  AND2X1 U67 ( .IN1(n52), .IN2(n7), .Q(n15) );
  AND2X1 U68 ( .IN1(n51), .IN2(n7), .Q(n14) );
  AND2X1 U69 ( .IN1(n50), .IN2(n7), .Q(n13) );
  AND2X1 U70 ( .IN1(n49), .IN2(n7), .Q(n12) );
  AND2X1 U71 ( .IN1(n48), .IN2(n7), .Q(n11) );
  AND2X1 U72 ( .IN1(n47), .IN2(n7), .Q(n10) );
  AO22X1 U73 ( .IN1(SH[5]), .IN2(n78), .IN3(n46), .IN4(n7), .Q(n9) );
  AND2X1 U78 ( .IN1(n115), .IN2(n44), .Q(n78) );
  AND2X1 U79 ( .IN1(n114), .IN2(n44), .Q(n77) );
  AND2X1 U80 ( .IN1(n113), .IN2(n44), .Q(n76) );
  AND2X1 U81 ( .IN1(n112), .IN2(n44), .Q(n75) );
  AND2X1 U82 ( .IN1(n111), .IN2(n44), .Q(n74) );
  AND2X1 U83 ( .IN1(n110), .IN2(n44), .Q(n73) );
  AND2X1 U84 ( .IN1(n109), .IN2(n44), .Q(n72) );
  AND2X1 U85 ( .IN1(n108), .IN2(n44), .Q(n71) );
  AND2X1 U86 ( .IN1(n107), .IN2(n44), .Q(n70) );
  AND2X1 U87 ( .IN1(n106), .IN2(n44), .Q(n69) );
  AND2X1 U88 ( .IN1(n105), .IN2(n44), .Q(n68) );
  AND2X1 U89 ( .IN1(n104), .IN2(n44), .Q(n67) );
  AND2X1 U90 ( .IN1(n103), .IN2(n44), .Q(n66) );
  AND2X1 U91 ( .IN1(n102), .IN2(n44), .Q(n65) );
  AND2X1 U92 ( .IN1(n101), .IN2(n44), .Q(n64) );
  AND2X1 U93 ( .IN1(n100), .IN2(n44), .Q(n63) );
  AO22X1 U94 ( .IN1(SH[4]), .IN2(n115), .IN3(n99), .IN4(n44), .Q(n62) );
  AO22X1 U95 ( .IN1(SH[4]), .IN2(n114), .IN3(n98), .IN4(n44), .Q(n61) );
  AO22X1 U96 ( .IN1(SH[4]), .IN2(n113), .IN3(n97), .IN4(n44), .Q(n60) );
  AO22X1 U97 ( .IN1(SH[4]), .IN2(n112), .IN3(n96), .IN4(n44), .Q(n59) );
  AO22X1 U98 ( .IN1(SH[4]), .IN2(n111), .IN3(n95), .IN4(n44), .Q(n58) );
  AO22X1 U99 ( .IN1(SH[4]), .IN2(n110), .IN3(n94), .IN4(n44), .Q(n57) );
  AO22X1 U100 ( .IN1(SH[4]), .IN2(n109), .IN3(n93), .IN4(n44), .Q(n56) );
  AO22X1 U101 ( .IN1(SH[4]), .IN2(n108), .IN3(n92), .IN4(n44), .Q(n55) );
  AO22X1 U102 ( .IN1(SH[4]), .IN2(n107), .IN3(n91), .IN4(n44), .Q(n54) );
  AO22X1 U103 ( .IN1(SH[4]), .IN2(n106), .IN3(n90), .IN4(n44), .Q(n53) );
  AO22X1 U104 ( .IN1(SH[4]), .IN2(n105), .IN3(n89), .IN4(n44), .Q(n52) );
  AO22X1 U105 ( .IN1(SH[4]), .IN2(n104), .IN3(n88), .IN4(n44), .Q(n51) );
  AO22X1 U106 ( .IN1(SH[4]), .IN2(n103), .IN3(n87), .IN4(n44), .Q(n50) );
  AO22X1 U107 ( .IN1(SH[4]), .IN2(n102), .IN3(n86), .IN4(n44), .Q(n49) );
  AO22X1 U108 ( .IN1(SH[4]), .IN2(n101), .IN3(n85), .IN4(n44), .Q(n48) );
  AO22X1 U109 ( .IN1(SH[4]), .IN2(n100), .IN3(n84), .IN4(n44), .Q(n47) );
  AO22X1 U110 ( .IN1(n44), .IN2(n83), .IN3(n99), .IN4(SH[4]), .Q(n46) );
  AND2X1 U115 ( .IN1(n152), .IN2(n81), .Q(n115) );
  AND2X1 U116 ( .IN1(n151), .IN2(n81), .Q(n114) );
  AND2X1 U117 ( .IN1(n150), .IN2(n81), .Q(n113) );
  AND2X1 U118 ( .IN1(n149), .IN2(n81), .Q(n112) );
  AND2X1 U119 ( .IN1(n148), .IN2(n81), .Q(n111) );
  AND2X1 U120 ( .IN1(n147), .IN2(n81), .Q(n110) );
  AND2X1 U121 ( .IN1(n146), .IN2(n81), .Q(n109) );
  AND2X1 U122 ( .IN1(n145), .IN2(n81), .Q(n108) );
  AO22X1 U123 ( .IN1(SH[3]), .IN2(n152), .IN3(n144), .IN4(n81), .Q(n107) );
  AO22X1 U124 ( .IN1(SH[3]), .IN2(n151), .IN3(n143), .IN4(n81), .Q(n106) );
  AO22X1 U125 ( .IN1(SH[3]), .IN2(n150), .IN3(n142), .IN4(n81), .Q(n105) );
  AO22X1 U126 ( .IN1(SH[3]), .IN2(n149), .IN3(n141), .IN4(n81), .Q(n104) );
  AO22X1 U127 ( .IN1(SH[3]), .IN2(n148), .IN3(n140), .IN4(n81), .Q(n103) );
  AO22X1 U128 ( .IN1(SH[3]), .IN2(n147), .IN3(n139), .IN4(n81), .Q(n102) );
  AO22X1 U129 ( .IN1(SH[3]), .IN2(n146), .IN3(n138), .IN4(n81), .Q(n101) );
  AO22X1 U130 ( .IN1(SH[3]), .IN2(n145), .IN3(n137), .IN4(n81), .Q(n100) );
  AO22X1 U131 ( .IN1(SH[3]), .IN2(n144), .IN3(n136), .IN4(n81), .Q(n99) );
  AO22X1 U132 ( .IN1(SH[3]), .IN2(n143), .IN3(n135), .IN4(n81), .Q(n98) );
  AO22X1 U133 ( .IN1(SH[3]), .IN2(n142), .IN3(n134), .IN4(n81), .Q(n97) );
  AO22X1 U134 ( .IN1(SH[3]), .IN2(n141), .IN3(n133), .IN4(n81), .Q(n96) );
  AO22X1 U135 ( .IN1(SH[3]), .IN2(n140), .IN3(n132), .IN4(n81), .Q(n95) );
  AO22X1 U136 ( .IN1(SH[3]), .IN2(n139), .IN3(n131), .IN4(n81), .Q(n94) );
  AO22X1 U137 ( .IN1(SH[3]), .IN2(n138), .IN3(n130), .IN4(n81), .Q(n93) );
  AO22X1 U138 ( .IN1(SH[3]), .IN2(n137), .IN3(n129), .IN4(n81), .Q(n92) );
  AO22X1 U139 ( .IN1(SH[3]), .IN2(n136), .IN3(n128), .IN4(n81), .Q(n91) );
  AO22X1 U140 ( .IN1(SH[3]), .IN2(n135), .IN3(n127), .IN4(n81), .Q(n90) );
  AO22X1 U141 ( .IN1(SH[3]), .IN2(n134), .IN3(n126), .IN4(n81), .Q(n89) );
  AO22X1 U142 ( .IN1(SH[3]), .IN2(n133), .IN3(n125), .IN4(n81), .Q(n88) );
  AO22X1 U143 ( .IN1(SH[3]), .IN2(n132), .IN3(n124), .IN4(n81), .Q(n87) );
  AO22X1 U144 ( .IN1(SH[3]), .IN2(n131), .IN3(n123), .IN4(n81), .Q(n86) );
  AO22X1 U145 ( .IN1(SH[3]), .IN2(n130), .IN3(n122), .IN4(n81), .Q(n85) );
  AO22X1 U146 ( .IN1(SH[3]), .IN2(n129), .IN3(n121), .IN4(n81), .Q(n84) );
  AO22X1 U147 ( .IN1(n81), .IN2(n120), .IN3(n128), .IN4(SH[3]), .Q(n83) );
  AND2X1 U152 ( .IN1(n189), .IN2(n118), .Q(n152) );
  AND2X1 U153 ( .IN1(n188), .IN2(n118), .Q(n151) );
  AND2X1 U154 ( .IN1(n187), .IN2(n118), .Q(n150) );
  AND2X1 U155 ( .IN1(n186), .IN2(n118), .Q(n149) );
  AO22X1 U156 ( .IN1(SH[2]), .IN2(n189), .IN3(n185), .IN4(n118), .Q(n148) );
  AO22X1 U157 ( .IN1(SH[2]), .IN2(n188), .IN3(n184), .IN4(n118), .Q(n147) );
  AO22X1 U158 ( .IN1(SH[2]), .IN2(n187), .IN3(n183), .IN4(n118), .Q(n146) );
  AO22X1 U159 ( .IN1(SH[2]), .IN2(n186), .IN3(n182), .IN4(n118), .Q(n145) );
  AO22X1 U160 ( .IN1(SH[2]), .IN2(n185), .IN3(n181), .IN4(n118), .Q(n144) );
  AO22X1 U161 ( .IN1(SH[2]), .IN2(n184), .IN3(n180), .IN4(n118), .Q(n143) );
  AO22X1 U162 ( .IN1(SH[2]), .IN2(n183), .IN3(n179), .IN4(n118), .Q(n142) );
  AO22X1 U163 ( .IN1(SH[2]), .IN2(n182), .IN3(n178), .IN4(n118), .Q(n141) );
  AO22X1 U164 ( .IN1(SH[2]), .IN2(n181), .IN3(n177), .IN4(n118), .Q(n140) );
  AO22X1 U165 ( .IN1(SH[2]), .IN2(n180), .IN3(n176), .IN4(n118), .Q(n139) );
  AO22X1 U166 ( .IN1(SH[2]), .IN2(n179), .IN3(n175), .IN4(n118), .Q(n138) );
  AO22X1 U167 ( .IN1(SH[2]), .IN2(n178), .IN3(n174), .IN4(n118), .Q(n137) );
  AO22X1 U168 ( .IN1(SH[2]), .IN2(n177), .IN3(n173), .IN4(n118), .Q(n136) );
  AO22X1 U169 ( .IN1(SH[2]), .IN2(n176), .IN3(n172), .IN4(n118), .Q(n135) );
  AO22X1 U170 ( .IN1(SH[2]), .IN2(n175), .IN3(n171), .IN4(n118), .Q(n134) );
  AO22X1 U171 ( .IN1(SH[2]), .IN2(n174), .IN3(n170), .IN4(n118), .Q(n133) );
  AO22X1 U172 ( .IN1(SH[2]), .IN2(n173), .IN3(n169), .IN4(n118), .Q(n132) );
  AO22X1 U173 ( .IN1(SH[2]), .IN2(n172), .IN3(n168), .IN4(n118), .Q(n131) );
  AO22X1 U174 ( .IN1(SH[2]), .IN2(n171), .IN3(n167), .IN4(n118), .Q(n130) );
  AO22X1 U175 ( .IN1(SH[2]), .IN2(n170), .IN3(n166), .IN4(n118), .Q(n129) );
  AO22X1 U176 ( .IN1(SH[2]), .IN2(n169), .IN3(n165), .IN4(n118), .Q(n128) );
  AO22X1 U177 ( .IN1(SH[2]), .IN2(n168), .IN3(n164), .IN4(n118), .Q(n127) );
  AO22X1 U178 ( .IN1(SH[2]), .IN2(n167), .IN3(n163), .IN4(n118), .Q(n126) );
  AO22X1 U179 ( .IN1(SH[2]), .IN2(n166), .IN3(n162), .IN4(n118), .Q(n125) );
  AO22X1 U180 ( .IN1(SH[2]), .IN2(n165), .IN3(n161), .IN4(n118), .Q(n124) );
  AO22X1 U181 ( .IN1(SH[2]), .IN2(n164), .IN3(n160), .IN4(n118), .Q(n123) );
  AO22X1 U182 ( .IN1(SH[2]), .IN2(n163), .IN3(n159), .IN4(n118), .Q(n122) );
  AO22X1 U183 ( .IN1(SH[2]), .IN2(n162), .IN3(n158), .IN4(n118), .Q(n121) );
  AO22X1 U184 ( .IN1(n118), .IN2(n157), .IN3(n161), .IN4(SH[2]), .Q(n120) );
  AND2X1 U189 ( .IN1(n225), .IN2(n155), .Q(n189) );
  AND2X1 U190 ( .IN1(n224), .IN2(n155), .Q(n188) );
  AO22X1 U191 ( .IN1(SH[1]), .IN2(n225), .IN3(n223), .IN4(n155), .Q(n187) );
  AO22X1 U192 ( .IN1(SH[1]), .IN2(n224), .IN3(n222), .IN4(n155), .Q(n186) );
  AO22X1 U193 ( .IN1(SH[1]), .IN2(n223), .IN3(n221), .IN4(n155), .Q(n185) );
  AO22X1 U194 ( .IN1(SH[1]), .IN2(n222), .IN3(n220), .IN4(n155), .Q(n184) );
  AO22X1 U195 ( .IN1(SH[1]), .IN2(n221), .IN3(n219), .IN4(n155), .Q(n183) );
  AO22X1 U196 ( .IN1(SH[1]), .IN2(n220), .IN3(n218), .IN4(n155), .Q(n182) );
  AO22X1 U197 ( .IN1(SH[1]), .IN2(n219), .IN3(n217), .IN4(n155), .Q(n181) );
  AO22X1 U198 ( .IN1(SH[1]), .IN2(n218), .IN3(n216), .IN4(n155), .Q(n180) );
  AO22X1 U199 ( .IN1(SH[1]), .IN2(n217), .IN3(n215), .IN4(n155), .Q(n179) );
  AO22X1 U200 ( .IN1(SH[1]), .IN2(n216), .IN3(n214), .IN4(n155), .Q(n178) );
  AO22X1 U201 ( .IN1(SH[1]), .IN2(n215), .IN3(n213), .IN4(n155), .Q(n177) );
  AO22X1 U202 ( .IN1(SH[1]), .IN2(n214), .IN3(n212), .IN4(n155), .Q(n176) );
  AO22X1 U203 ( .IN1(SH[1]), .IN2(n213), .IN3(n211), .IN4(n155), .Q(n175) );
  AO22X1 U204 ( .IN1(SH[1]), .IN2(n212), .IN3(n210), .IN4(n155), .Q(n174) );
  AO22X1 U205 ( .IN1(SH[1]), .IN2(n211), .IN3(n209), .IN4(n155), .Q(n173) );
  AO22X1 U206 ( .IN1(SH[1]), .IN2(n210), .IN3(n208), .IN4(n155), .Q(n172) );
  AO22X1 U207 ( .IN1(SH[1]), .IN2(n209), .IN3(n207), .IN4(n155), .Q(n171) );
  AO22X1 U208 ( .IN1(SH[1]), .IN2(n208), .IN3(n206), .IN4(n155), .Q(n170) );
  AO22X1 U209 ( .IN1(SH[1]), .IN2(n207), .IN3(n205), .IN4(n155), .Q(n169) );
  AO22X1 U210 ( .IN1(SH[1]), .IN2(n206), .IN3(n204), .IN4(n155), .Q(n168) );
  AO22X1 U211 ( .IN1(SH[1]), .IN2(n205), .IN3(n203), .IN4(n155), .Q(n167) );
  AO22X1 U212 ( .IN1(SH[1]), .IN2(n204), .IN3(n202), .IN4(n155), .Q(n166) );
  AO22X1 U213 ( .IN1(SH[1]), .IN2(n203), .IN3(n201), .IN4(n155), .Q(n165) );
  AO22X1 U214 ( .IN1(SH[1]), .IN2(n202), .IN3(n200), .IN4(n155), .Q(n164) );
  AO22X1 U215 ( .IN1(SH[1]), .IN2(n201), .IN3(n199), .IN4(n155), .Q(n163) );
  AO22X1 U216 ( .IN1(SH[1]), .IN2(n200), .IN3(n198), .IN4(n155), .Q(n162) );
  AO22X1 U217 ( .IN1(SH[1]), .IN2(n199), .IN3(n197), .IN4(n155), .Q(n161) );
  AO22X1 U218 ( .IN1(SH[1]), .IN2(n198), .IN3(n196), .IN4(n155), .Q(n160) );
  AO22X1 U219 ( .IN1(SH[1]), .IN2(n197), .IN3(n195), .IN4(n155), .Q(n159) );
  AO22X1 U220 ( .IN1(SH[1]), .IN2(n196), .IN3(n194), .IN4(n155), .Q(n158) );
  AO22X1 U221 ( .IN1(n193), .IN2(n155), .IN3(n195), .IN4(SH[1]), .Q(n157) );
  AND2X1 U225 ( .IN1(n191), .IN2(A[32]), .Q(n225) );
  AO22X1 U226 ( .IN1(A[32]), .IN2(SH[0]), .IN3(n191), .IN4(A[31]), .Q(n224) );
  AO22X1 U227 ( .IN1(A[31]), .IN2(SH[0]), .IN3(n191), .IN4(A[30]), .Q(n223) );
  AO22X1 U228 ( .IN1(A[30]), .IN2(SH[0]), .IN3(n191), .IN4(A[29]), .Q(n222) );
  AO22X1 U229 ( .IN1(A[29]), .IN2(SH[0]), .IN3(n191), .IN4(A[28]), .Q(n221) );
  AO22X1 U230 ( .IN1(A[28]), .IN2(SH[0]), .IN3(n191), .IN4(A[27]), .Q(n220) );
  AO22X1 U231 ( .IN1(A[27]), .IN2(SH[0]), .IN3(n191), .IN4(A[26]), .Q(n219) );
  AO22X1 U232 ( .IN1(A[26]), .IN2(SH[0]), .IN3(n191), .IN4(A[25]), .Q(n218) );
  AO22X1 U233 ( .IN1(A[25]), .IN2(SH[0]), .IN3(n191), .IN4(A[24]), .Q(n217) );
  AO22X1 U234 ( .IN1(A[24]), .IN2(SH[0]), .IN3(n191), .IN4(A[23]), .Q(n216) );
  AO22X1 U235 ( .IN1(A[23]), .IN2(SH[0]), .IN3(n191), .IN4(A[22]), .Q(n215) );
  AO22X1 U236 ( .IN1(A[22]), .IN2(SH[0]), .IN3(n191), .IN4(A[21]), .Q(n214) );
  AO22X1 U237 ( .IN1(A[21]), .IN2(SH[0]), .IN3(n191), .IN4(A[20]), .Q(n213) );
  AO22X1 U238 ( .IN1(A[20]), .IN2(SH[0]), .IN3(n191), .IN4(A[19]), .Q(n212) );
  AO22X1 U239 ( .IN1(A[19]), .IN2(SH[0]), .IN3(n191), .IN4(A[18]), .Q(n211) );
  AO22X1 U240 ( .IN1(A[18]), .IN2(SH[0]), .IN3(n191), .IN4(A[17]), .Q(n210) );
  AO22X1 U241 ( .IN1(A[17]), .IN2(SH[0]), .IN3(n191), .IN4(A[16]), .Q(n209) );
  AO22X1 U242 ( .IN1(A[16]), .IN2(SH[0]), .IN3(n191), .IN4(A[15]), .Q(n208) );
  AO22X1 U243 ( .IN1(A[15]), .IN2(SH[0]), .IN3(n191), .IN4(A[14]), .Q(n207) );
  AO22X1 U244 ( .IN1(A[14]), .IN2(SH[0]), .IN3(n191), .IN4(A[13]), .Q(n206) );
  AO22X1 U245 ( .IN1(A[13]), .IN2(SH[0]), .IN3(n191), .IN4(A[12]), .Q(n205) );
  AO22X1 U246 ( .IN1(A[12]), .IN2(SH[0]), .IN3(n191), .IN4(A[11]), .Q(n204) );
  AO22X1 U247 ( .IN1(A[11]), .IN2(SH[0]), .IN3(n191), .IN4(A[10]), .Q(n203) );
  AO22X1 U248 ( .IN1(A[10]), .IN2(SH[0]), .IN3(n191), .IN4(A[9]), .Q(n202) );
  AO22X1 U249 ( .IN1(A[9]), .IN2(SH[0]), .IN3(n191), .IN4(A[8]), .Q(n201) );
  AO22X1 U250 ( .IN1(A[8]), .IN2(SH[0]), .IN3(n191), .IN4(A[7]), .Q(n200) );
  AO22X1 U251 ( .IN1(A[7]), .IN2(SH[0]), .IN3(n191), .IN4(A[6]), .Q(n199) );
  AO22X1 U252 ( .IN1(A[6]), .IN2(SH[0]), .IN3(n191), .IN4(A[5]), .Q(n198) );
  AO22X1 U253 ( .IN1(A[5]), .IN2(SH[0]), .IN3(n191), .IN4(A[4]), .Q(n197) );
  AO22X1 U254 ( .IN1(A[4]), .IN2(SH[0]), .IN3(n191), .IN4(A[3]), .Q(n196) );
  AO22X1 U255 ( .IN1(A[3]), .IN2(SH[0]), .IN3(n191), .IN4(A[2]), .Q(n195) );
  AO22X1 U256 ( .IN1(A[2]), .IN2(SH[0]), .IN3(n191), .IN4(A[1]), .Q(n194) );
  AND2X1 U257 ( .IN1(SH[0]), .IN2(A[1]), .Q(n193) );
  INVX0 U263 ( .INP(SH[1]), .ZN(n155) );
  INVX0 U264 ( .INP(SH[0]), .ZN(n191) );
  INVX0 U265 ( .INP(SH[2]), .ZN(n118) );
  INVX0 U266 ( .INP(SH[3]), .ZN(n81) );
  INVX0 U267 ( .INP(SH[4]), .ZN(n44) );
  INVX0 U268 ( .INP(SH[5]), .ZN(n7) );
  NOR2X0 U269 ( .IN1(SH[7]), .IN2(SH[6]), .QN(n307) );
endmodule


module thumb ( read_instruction_n, instruction_address, instruction, 
        read_data_n, write_data_n, data_address, data, reset_n, clk );
  output [31:0] instruction_address;
  input [15:0] instruction;
  output [31:0] data_address;
  inout [31:0] data;
  input reset_n, clk;
  output read_instruction_n, read_data_n, write_data_n;
  wire   N136, N307, N308, N310, N311, N313, N315, N318, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N435, N436, N437, N438,
         N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, \R[7][31] , \R[7][30] ,
         \R[7][29] , \R[7][28] , \R[7][27] , \R[7][26] , \R[7][25] ,
         \R[7][24] , \R[7][23] , \R[7][22] , \R[7][21] , \R[7][20] ,
         \R[7][19] , \R[7][18] , \R[7][17] , \R[7][16] , \R[7][15] ,
         \R[7][14] , \R[7][13] , \R[7][12] , \R[7][11] , \R[7][10] , \R[7][9] ,
         \R[7][8] , \R[7][7] , \R[7][6] , \R[7][5] , \R[7][4] , \R[7][3] ,
         \R[7][2] , \R[7][1] , \R[7][0] , \R[6][31] , \R[6][30] , \R[6][29] ,
         \R[6][28] , \R[6][27] , \R[6][26] , \R[6][25] , \R[6][24] ,
         \R[6][23] , \R[6][22] , \R[6][21] , \R[6][20] , \R[6][19] ,
         \R[6][18] , \R[6][17] , \R[6][16] , \R[6][15] , \R[6][14] ,
         \R[6][13] , \R[6][12] , \R[6][11] , \R[6][10] , \R[6][9] , \R[6][8] ,
         \R[6][7] , \R[6][6] , \R[6][5] , \R[6][4] , \R[6][3] , \R[6][2] ,
         \R[6][1] , \R[6][0] , \R[5][31] , \R[5][30] , \R[5][29] , \R[5][28] ,
         \R[5][27] , \R[5][26] , \R[5][25] , \R[5][24] , \R[5][23] ,
         \R[5][22] , \R[5][21] , \R[5][20] , \R[5][19] , \R[5][18] ,
         \R[5][17] , \R[5][16] , \R[5][15] , \R[5][14] , \R[5][13] ,
         \R[5][12] , \R[5][11] , \R[5][10] , \R[5][9] , \R[5][8] , \R[5][7] ,
         \R[5][6] , \R[5][5] , \R[5][4] , \R[5][3] , \R[5][2] , \R[5][1] ,
         \R[5][0] , \R[4][31] , \R[4][30] , \R[4][29] , \R[4][28] , \R[4][27] ,
         \R[4][26] , \R[4][25] , \R[4][24] , \R[4][23] , \R[4][22] ,
         \R[4][21] , \R[4][20] , \R[4][19] , \R[4][18] , \R[4][17] ,
         \R[4][16] , \R[4][15] , \R[4][14] , \R[4][13] , \R[4][12] ,
         \R[4][11] , \R[4][10] , \R[4][9] , \R[4][8] , \R[4][7] , \R[4][6] ,
         \R[4][5] , \R[4][4] , \R[4][3] , \R[4][2] , \R[4][1] , \R[4][0] ,
         \R[3][31] , \R[3][30] , \R[3][29] , \R[3][28] , \R[3][27] ,
         \R[3][26] , \R[3][25] , \R[3][24] , \R[3][23] , \R[3][22] ,
         \R[3][21] , \R[3][20] , \R[3][19] , \R[3][18] , \R[3][17] ,
         \R[3][16] , \R[3][15] , \R[3][14] , \R[3][13] , \R[3][12] ,
         \R[3][11] , \R[3][10] , \R[3][9] , \R[3][8] , \R[3][7] , \R[3][6] ,
         \R[3][5] , \R[3][4] , \R[3][3] , \R[3][2] , \R[3][1] , \R[3][0] ,
         \R[2][31] , \R[2][30] , \R[2][29] , \R[2][28] , \R[2][27] ,
         \R[2][26] , \R[2][25] , \R[2][24] , \R[2][23] , \R[2][22] ,
         \R[2][21] , \R[2][20] , \R[2][19] , \R[2][18] , \R[2][17] ,
         \R[2][16] , \R[2][15] , \R[2][14] , \R[2][13] , \R[2][12] ,
         \R[2][11] , \R[2][10] , \R[2][9] , \R[2][8] , \R[2][7] , \R[2][6] ,
         \R[2][5] , \R[2][4] , \R[2][3] , \R[2][2] , \R[2][1] , \R[2][0] ,
         \R[1][31] , \R[1][30] , \R[1][29] , \R[1][28] , \R[1][27] ,
         \R[1][26] , \R[1][25] , \R[1][24] , \R[1][23] , \R[1][22] ,
         \R[1][21] , \R[1][20] , \R[1][19] , \R[1][18] , \R[1][17] ,
         \R[1][16] , \R[1][15] , \R[1][14] , \R[1][13] , \R[1][12] ,
         \R[1][11] , \R[1][10] , \R[1][9] , \R[1][8] , \R[1][7] , \R[1][6] ,
         \R[1][5] , \R[1][4] , \R[1][3] , \R[1][2] , \R[1][1] , \R[1][0] ,
         \R[0][31] , \R[0][30] , \R[0][29] , \R[0][28] , \R[0][27] ,
         \R[0][26] , \R[0][25] , \R[0][24] , \R[0][23] , \R[0][22] ,
         \R[0][21] , \R[0][20] , \R[0][19] , \R[0][18] , \R[0][17] ,
         \R[0][16] , \R[0][15] , \R[0][14] , \R[0][13] , \R[0][12] ,
         \R[0][11] , \R[0][10] , \R[0][9] , \R[0][8] , \R[0][7] , \R[0][6] ,
         \R[0][5] , \R[0][4] , \R[0][3] , \R[0][2] , \R[0][1] , \R[0][0] ,
         N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477,
         N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488,
         N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499,
         N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510,
         N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521,
         N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532,
         N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543,
         N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554,
         N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565,
         N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576,
         N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587,
         N588, N589, N590, N591, N592, N593, N594, N1187, N1188, N1189, N1190,
         N1191, N1192, N1254, N1255, N1735, N1736, N1737, N1738, N1739, N1740,
         N1741, N1742, N1743, N1744, N1745, N1746, N1747, N1748, N1749, N1750,
         N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, N1759, N1760,
         N1761, N1762, N1763, N1764, N1765, N1766, N1767, N1770, N1771, N1772,
         N1773, N1774, N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782,
         N1783, N1784, N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792,
         N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802,
         N1803, N1804, N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812,
         N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822,
         N1823, N1824, N1825, N1826, N1827, N1828, N1829, N1830, N1831, N1864,
         N1865, N1866, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874,
         N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884,
         N1885, N1886, N1887, N1888, N1889, N1890, N1891, N1892, N1893, N1894,
         N1895, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993,
         N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003,
         N3004, N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013,
         N3014, N3015, N3016, N4110, N4111, N4112, N4113, N4114, N4115, N4116,
         N4117, N4118, N4119, N4120, N4121, N4122, N4123, N4124, N4125, N4126,
         N4127, N4128, N4129, N4130, N4131, N4132, N4133, N4134, N4135, N4136,
         N4137, N4138, N4139, N4140, N4141, N4351, N4352, N4353, N4354, N4355,
         N4356, N4357, N4358, N4359, N4360, N4361, N4362, N4363, N4364, N4365,
         N4366, N4367, N4368, N4369, N4370, N4371, N4372, N4373, N4374, N4375,
         N4376, N4377, N4378, N4379, N4380, N4381, N4382, N4481, N4482, N4483,
         N4484, N4485, N4486, N4487, N4488, N4489, N4490, N4491, N4492, N4493,
         N4494, N4495, N4496, N4497, N4498, N4499, N4500, N4501, N4502, N4503,
         N4504, N4505, N4506, N4507, N4508, N4509, N4510, N4511, N4512, N4513,
         N4514, N4515, N4516, N4517, N4518, N4519, N4520, N4521, N4522, N4523,
         N4524, N4525, N4526, N4527, N4528, N4529, N4530, N4531, N4532, N4533,
         N4534, N4535, N4536, N4537, N4538, N4539, N4540, N4541, N4542, N4543,
         N4544, N4545, N4546, N4547, N4548, N4549, N4550, N4551, N4552, N4553,
         N4554, N4555, N4556, N4557, N4558, N4559, N4560, N4561, N4562, N4563,
         N4564, N4565, N4566, N4567, N4568, N4569, N4570, N4571, N4572, N4573,
         N4574, N4575, N4576, N4577, N4578, N4579, N4580, N4581, N4582, N4583,
         N4584, N4585, N4586, N4587, N4588, N4589, N4590, N4591, N4592, N4593,
         N4594, N4595, N4596, N4597, N4598, N4599, N4600, N4601, N4602, N4603,
         N4604, N4605, N4606, N4607, N4608, N4609, N4610, N4611, N4677, N4710,
         N4711, N4712, N4713, N4714, N4715, N4716, N4717, N4718, N4719, N4720,
         N4721, N4722, N4723, N4724, N4725, N4726, N4727, N4728, N4729, N4730,
         N4731, N4732, N4733, N4734, N4735, N4736, N4737, N4738, N4739, N4740,
         N4741, N4742, N4743, N4744, N4745, N4746, N4747, N4748, N4749, N4750,
         N4751, N4752, N4753, N4754, N4755, N4756, N4757, N4758, N4759, N4760,
         N4761, N4762, N4763, N4764, N4765, N4766, N4767, N4768, N4769, N4770,
         N4771, N4772, N4773, N4774, N4775, N4776, N4777, N4778, N4779, N4780,
         N4781, N4782, N4783, N4784, N4785, N4786, N4787, N4788, N4789, N4790,
         N4791, N4792, N4793, N4794, N4795, N4796, N4797, N4798, N4799, N4800,
         N4801, N4802, N4803, N4804, N4805, N4806, N4807, N4808, N4809, N4813,
         N4814, N4815, N4816, N4817, N4818, N4819, N4820, N4821, N4822, N4823,
         N4824, N4825, N4826, N4827, N4828, N4829, N4830, N4831, N4832, N4833,
         N4834, N4835, N4836, N4837, N4838, N4839, N4840, N4841, N4842, N4843,
         N4844, N4845, N4846, N4847, N4848, N4849, N4850, N4851, N4852, N4853,
         N4854, N4855, N4856, N4857, N4858, N4859, N4860, N4861, N4862, N4863,
         N4864, N4865, N4866, N4867, N4868, N4869, N4870, N4871, N4872, N4873,
         N4874, N4875, N4876, N4877, N4879, N4880, N4881, N4882, N4883, N4884,
         N4885, N4886, N4887, N4888, N4889, N4890, N4891, N4892, N4893, N4894,
         N4895, N4896, N4897, N4898, N4899, N4900, N4901, N4902, N4903, N4904,
         N4905, N4906, N4907, N4908, N4909, N4910, N4911, N4915, N4916, N4917,
         N4918, N4919, N4920, N4921, N4922, N4923, N4924, N4925, N4926, N4927,
         N4928, N4929, N4930, N4931, N4932, N4933, N4934, N4935, N4936, N4937,
         N4938, N4939, N4940, N4941, N4942, N4943, N4944, N4945, N4946, N4947,
         N4948, N4949, N4950, N4951, N4952, N4953, N4954, N4955, N4956, N4957,
         N4958, N4959, N4960, N4961, N4962, N4963, N4964, N4965, N4966, N4967,
         N4968, N4969, N4970, N4971, N4972, N4973, N4974, N4975, N4976, N4977,
         N4978, N4979, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N4988,
         N4989, N4990, N4991, N4992, N4993, N4994, N4995, N4996, N4997, N4998,
         N4999, N5000, N5001, N5002, N5003, N5004, N5005, N5006, N5007, N5008,
         N5009, N5010, N5011, N5012, N5046, N5047, N5048, N5049, N5050, N5051,
         N5052, N5053, N5054, N5055, N5056, N5057, N5058, N5059, N5060, N5061,
         N5062, N5063, N5064, N5065, N5066, N5067, N5068, N5069, N5070, N5071,
         N5072, N5073, N5074, N5075, N5076, N5077, N5162, N5163, N5164, N5165,
         N5166, N5167, N5168, N5169, N5170, N5171, N5172, N5173, N5174, N5175,
         N5176, N5177, N5178, N5179, N5180, N5181, N5182, N5183, N5184, N5185,
         N5186, N5187, N5188, N5189, N5190, N5191, N5192, N5193, N5194, N5195,
         N5196, N5197, N5198, N5199, N5200, N5201, N5202, N5203, N5204, N5205,
         N5206, N5207, N5208, N5209, N5210, N5211, N5212, N5213, N5214, N5215,
         N5216, N5217, N5218, N5219, N5220, N5221, N5222, N5223, N5224, N5225,
         N5226, N5260, N5261, N5262, N5263, N5264, N5265, N5266, N5267, N5268,
         N5269, N5270, N5271, N5272, N5273, N5274, N5275, N5276, N5277, N5278,
         N5279, N5280, N5281, N5282, N5283, N5284, N5285, N5286, N5287, N5288,
         N5289, N5290, N5291, N5292, N5622, N5623, N5624, N5625, N5626, N5627,
         N5628, N5629, N5630, N5631, N5632, N5633, N5634, N5635, N5636, N5637,
         N5638, N5639, N5640, N5641, N5642, N5643, N5644, N5645, N5646, N5647,
         N5648, N5649, N5650, N5651, N5652, N5653, N6323, N6325, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, \U3/U85/Z_4 ,
         \U3/U87/Z_0 , \U3/U87/Z_1 , \U3/U87/Z_2 , \U3/U87/Z_3 , \U3/U87/Z_4 ,
         \U3/U87/Z_5 , \U3/U87/Z_6 , \U3/U87/Z_7 , \U3/U87/Z_8 , \U3/U87/Z_9 ,
         \U3/U87/Z_10 , \U3/U87/Z_11 , \U3/U87/Z_12 , \U3/U87/Z_13 ,
         \U3/U87/Z_14 , \U3/U87/Z_15 , \U3/U87/Z_16 , \U3/U87/Z_17 ,
         \U3/U87/Z_18 , \U3/U87/Z_19 , \U3/U87/Z_20 , \U3/U87/Z_21 ,
         \U3/U87/Z_22 , \U3/U87/Z_23 , \U3/U87/Z_24 , \U3/U87/Z_25 ,
         \U3/U87/Z_26 , \U3/U87/Z_27 , \U3/U87/Z_28 , \U3/U87/Z_29 ,
         \U3/U87/Z_30 , \U3/U87/Z_31 , \U3/U88/Z_0 , \U3/U88/Z_1 ,
         \U3/U88/Z_2 , \U3/U88/Z_3 , \U3/U88/Z_4 , \U3/U88/Z_5 , \U3/U88/Z_6 ,
         \U3/U88/Z_7 , \U3/U88/Z_8 , \U3/U88/Z_9 , \U3/U88/Z_10 ,
         \U3/U88/Z_11 , \U3/U88/Z_12 , \U3/U88/Z_13 , \U3/U88/Z_14 ,
         \U3/U88/Z_15 , \U3/U88/Z_16 , \U3/U88/Z_17 , \U3/U88/Z_18 ,
         \U3/U88/Z_19 , \U3/U88/Z_20 , \U3/U88/Z_21 , \U3/U88/Z_22 ,
         \U3/U88/Z_23 , \U3/U88/Z_24 , \U3/U88/Z_25 , \U3/U88/Z_26 ,
         \U3/U88/Z_27 , \U3/U88/Z_28 , \U3/U88/Z_29 , \U3/U88/Z_30 ,
         \U3/U88/Z_31 , \U3/U88/Z_32 , \U3/U89/Z_0 , \U3/U90/Z_0 ,
         \U3/U91/Z_0 , \U3/U91/Z_1 , \U3/U91/Z_2 , \U3/U91/Z_3 , \U3/U91/Z_4 ,
         \U3/U91/Z_5 , \U3/U91/Z_6 , \U3/U91/Z_7 , \U3/U91/Z_8 , \U3/U91/Z_9 ,
         \U3/U91/Z_10 , \U3/U91/Z_11 , \U3/U91/Z_12 , \U3/U91/Z_13 ,
         \U3/U91/Z_14 , \U3/U91/Z_15 , \U3/U91/Z_16 , \U3/U91/Z_17 ,
         \U3/U91/Z_18 , \U3/U91/Z_19 , \U3/U91/Z_20 , \U3/U91/Z_21 ,
         \U3/U91/Z_22 , \U3/U91/Z_23 , \U3/U91/Z_24 , \U3/U91/Z_25 ,
         \U3/U91/Z_26 , \U3/U91/Z_27 , \U3/U91/Z_28 , \U3/U91/Z_29 ,
         \U3/U91/Z_30 , \U3/U91/Z_31 , \U3/U92/Z_0 , \U3/U92/Z_1 ,
         \U3/U92/Z_2 , \U3/U92/Z_3 , \U3/U92/Z_4 , \U3/U92/Z_5 , \U3/U92/Z_6 ,
         \U3/U92/Z_7 , \U3/U92/Z_8 , \U3/U92/Z_9 , \U3/U92/Z_10 ,
         \U3/U92/Z_11 , \U3/U93/Z_0 , n3573, n3574, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3700, n3704,
         n3705, n3711, n3713, n3714, n3715, n3716, n3719, n3720, n3721, n3723,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, \r1720/A[3] ,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230;
  wire   [31:0] IF_PC;
  wire   [5:0] ID_opcode;
  wire   [10:0] ID_imm_offset;
  wire   [31:0] ID_Rn;
  wire   [31:0] ID_Rd;
  wire   [31:0] ID_Rm_Rs;
  wire   [31:0] ID_PC;
  wire   [31:0] SP;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;
  assign read_instruction_n = 1'b0;

  DFFX1 \ID_opcode_reg[4]  ( .D(N1191), .CLK(clk), .Q(ID_opcode[4]), .QN(n3720) );
  DFFX1 \ID_opcode_reg[0]  ( .D(N1187), .CLK(clk), .Q(\U3/U85/Z_4 ), .QN(
        \r1720/A[3] ) );
  DFFX1 \ID_opcode_reg[1]  ( .D(N1188), .CLK(clk), .Q(n5695), .QN(n3723) );
  DFFX1 \ID_opcode_reg[2]  ( .D(N1189), .CLK(clk), .Q(ID_opcode[2]), .QN(n3716) );
  DFFX1 \ID_opcode_reg[3]  ( .D(N1190), .CLK(clk), .Q(ID_opcode[3]), .QN(n3719) );
  DFFX1 \ID_opcode_reg[5]  ( .D(N1192), .CLK(clk), .Q(n5696), .QN(n3721) );
  DFFASX1 write_data_n_reg ( .D(N6325), .CLK(clk), .SETB(reset_n), .Q(
        write_data_n), .QN(n9198) );
  DFFASX1 read_data_n_reg ( .D(N6323), .CLK(clk), .SETB(reset_n), .Q(
        read_data_n) );
  DFFX1 \ID_PC_reg[31]  ( .D(IF_PC[31]), .CLK(clk), .Q(ID_PC[31]) );
  DFFARX1 \PC_reg[31]  ( .D(N466), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[31]) );
  DFFX1 \ID_PC_reg[0]  ( .D(IF_PC[0]), .CLK(clk), .Q(n9172) );
  DFFARX1 \PC_reg[0]  ( .D(N435), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[0]) );
  DFFX1 \ID_PC_reg[1]  ( .D(IF_PC[1]), .CLK(clk), .Q(n9171) );
  DFFARX1 \PC_reg[1]  ( .D(N436), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[1]) );
  DFFX1 \ID_PC_reg[2]  ( .D(IF_PC[2]), .CLK(clk), .Q(ID_PC[2]) );
  DFFARX1 \PC_reg[2]  ( .D(N437), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[2]) );
  DFFX1 \ID_PC_reg[3]  ( .D(IF_PC[3]), .CLK(clk), .Q(ID_PC[3]) );
  DFFARX1 \PC_reg[3]  ( .D(N438), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[3]) );
  DFFX1 \ID_PC_reg[4]  ( .D(IF_PC[4]), .CLK(clk), .Q(ID_PC[4]) );
  DFFARX1 \PC_reg[4]  ( .D(N439), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[4]) );
  DFFX1 \ID_PC_reg[5]  ( .D(IF_PC[5]), .CLK(clk), .Q(ID_PC[5]) );
  DFFARX1 \PC_reg[5]  ( .D(N440), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[5]) );
  DFFX1 \ID_PC_reg[6]  ( .D(IF_PC[6]), .CLK(clk), .Q(ID_PC[6]) );
  DFFARX1 \PC_reg[6]  ( .D(N441), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[6]) );
  DFFX1 \ID_PC_reg[7]  ( .D(IF_PC[7]), .CLK(clk), .Q(ID_PC[7]) );
  DFFARX1 \PC_reg[7]  ( .D(N442), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[7]) );
  DFFX1 \ID_PC_reg[8]  ( .D(IF_PC[8]), .CLK(clk), .Q(ID_PC[8]) );
  DFFARX1 \PC_reg[8]  ( .D(N443), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[8]) );
  DFFX1 \ID_PC_reg[9]  ( .D(IF_PC[9]), .CLK(clk), .Q(ID_PC[9]) );
  DFFARX1 \PC_reg[9]  ( .D(N444), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[9]) );
  DFFX1 \ID_PC_reg[10]  ( .D(IF_PC[10]), .CLK(clk), .Q(ID_PC[10]) );
  DFFARX1 \PC_reg[10]  ( .D(N445), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[10]) );
  DFFX1 \ID_PC_reg[11]  ( .D(IF_PC[11]), .CLK(clk), .Q(ID_PC[11]) );
  DFFARX1 \PC_reg[11]  ( .D(N446), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[11]) );
  DFFX1 \ID_PC_reg[12]  ( .D(IF_PC[12]), .CLK(clk), .Q(ID_PC[12]) );
  DFFARX1 \PC_reg[12]  ( .D(N447), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[12]) );
  DFFX1 \ID_PC_reg[13]  ( .D(IF_PC[13]), .CLK(clk), .Q(ID_PC[13]) );
  DFFARX1 \PC_reg[13]  ( .D(N448), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[13]) );
  DFFX1 \ID_PC_reg[14]  ( .D(IF_PC[14]), .CLK(clk), .Q(ID_PC[14]) );
  DFFARX1 \PC_reg[14]  ( .D(N449), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[14]) );
  DFFX1 \ID_PC_reg[15]  ( .D(IF_PC[15]), .CLK(clk), .Q(ID_PC[15]) );
  DFFARX1 \PC_reg[15]  ( .D(N450), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[15]) );
  DFFX1 \ID_PC_reg[16]  ( .D(IF_PC[16]), .CLK(clk), .Q(ID_PC[16]) );
  DFFARX1 \PC_reg[16]  ( .D(N451), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[16]) );
  DFFX1 \ID_PC_reg[17]  ( .D(IF_PC[17]), .CLK(clk), .Q(ID_PC[17]) );
  DFFARX1 \PC_reg[17]  ( .D(N452), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[17]) );
  DFFX1 \ID_PC_reg[18]  ( .D(IF_PC[18]), .CLK(clk), .Q(ID_PC[18]) );
  DFFARX1 \PC_reg[18]  ( .D(N453), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[18]) );
  DFFX1 \ID_PC_reg[19]  ( .D(IF_PC[19]), .CLK(clk), .Q(ID_PC[19]) );
  DFFARX1 \PC_reg[19]  ( .D(N454), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[19]) );
  DFFX1 \ID_PC_reg[20]  ( .D(IF_PC[20]), .CLK(clk), .Q(ID_PC[20]) );
  DFFARX1 \PC_reg[20]  ( .D(N455), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[20]) );
  DFFX1 \ID_PC_reg[21]  ( .D(IF_PC[21]), .CLK(clk), .Q(ID_PC[21]) );
  DFFARX1 \PC_reg[21]  ( .D(N456), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[21]) );
  DFFX1 \ID_PC_reg[22]  ( .D(IF_PC[22]), .CLK(clk), .Q(ID_PC[22]) );
  DFFARX1 \PC_reg[22]  ( .D(N457), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[22]) );
  DFFX1 \ID_PC_reg[23]  ( .D(IF_PC[23]), .CLK(clk), .Q(ID_PC[23]) );
  DFFARX1 \PC_reg[23]  ( .D(N458), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[23]) );
  DFFX1 \ID_PC_reg[24]  ( .D(IF_PC[24]), .CLK(clk), .Q(ID_PC[24]) );
  DFFARX1 \PC_reg[24]  ( .D(N459), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[24]) );
  DFFX1 \ID_PC_reg[25]  ( .D(IF_PC[25]), .CLK(clk), .Q(ID_PC[25]) );
  DFFARX1 \PC_reg[25]  ( .D(N460), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[25]) );
  DFFX1 \ID_PC_reg[26]  ( .D(IF_PC[26]), .CLK(clk), .Q(ID_PC[26]) );
  DFFARX1 \PC_reg[26]  ( .D(N461), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[26]) );
  DFFX1 \ID_PC_reg[27]  ( .D(IF_PC[27]), .CLK(clk), .Q(ID_PC[27]) );
  DFFARX1 \PC_reg[27]  ( .D(N462), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[27]) );
  DFFX1 \ID_PC_reg[28]  ( .D(IF_PC[28]), .CLK(clk), .Q(ID_PC[28]) );
  DFFARX1 \PC_reg[28]  ( .D(N463), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[28]) );
  DFFX1 \ID_PC_reg[29]  ( .D(IF_PC[29]), .CLK(clk), .Q(ID_PC[29]) );
  DFFARX1 \PC_reg[29]  ( .D(N464), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[29]) );
  DFFX1 \ID_PC_reg[30]  ( .D(IF_PC[30]), .CLK(clk), .Q(ID_PC[30]) );
  DFFARX1 \PC_reg[30]  ( .D(N465), .CLK(clk), .RSTB(reset_n), .Q(
        instruction_address[30]) );
  DFFX1 \LR_reg[0]  ( .D(n4421), .CLK(clk), .Q(n9170) );
  DFFX1 V_Flag_reg ( .D(n4420), .CLK(clk), .Q(n9169) );
  DFFARX1 branch_taken_reg ( .D(n4419), .CLK(clk), .RSTB(reset_n), .Q(n9191), 
        .QN(n5701) );
  DFFX1 \IF_IR_reg[9]  ( .D(n4418), .CLK(clk), .Q(N136), .QN(n3711) );
  DFFX1 \IF_IR_reg[10]  ( .D(n4417), .CLK(clk), .Q(N315), .QN(n4422) );
  DFFX1 \IF_IR_reg[11]  ( .D(n4416), .CLK(clk), .Q(n9186), .QN(n5702) );
  DFFX1 \IF_IR_reg[12]  ( .D(n4415), .CLK(clk), .Q(n9187), .QN(n5689) );
  DFFX1 \IF_IR_reg[14]  ( .D(n4414), .CLK(clk), .Q(n9188), .QN(n5692) );
  DFFX1 \IF_IR_reg[15]  ( .D(n4413), .CLK(clk), .Q(n9185), .QN(n5705) );
  DFFX1 \IF_IR_reg[13]  ( .D(n4412), .CLK(clk), .Q(n9189), .QN(n5686) );
  DFFX1 \ID_imm_offset_reg[9]  ( .D(n4411), .CLK(clk), .Q(ID_imm_offset[9]), 
        .QN(n3705) );
  DFFX1 \ID_imm_offset_reg[10]  ( .D(n4410), .CLK(clk), .Q(ID_imm_offset[10]), 
        .QN(n3704) );
  DFFX1 \ID_cond_reg[1]  ( .D(n4409), .CLK(clk), .Q(n9168) );
  DFFX1 \ID_cond_reg[2]  ( .D(n4408), .CLK(clk), .Q(n9190) );
  DFFX1 \ID_cond_reg[3]  ( .D(n4407), .CLK(clk), .Q(n9167) );
  DFFX1 \IF_IR_reg[8]  ( .D(n4406), .CLK(clk), .Q(n5697), .QN(n3700) );
  DFFX1 \ID_cond_reg[0]  ( .D(n4405), .CLK(clk), .Q(n9166) );
  DFFX1 \ID_imm_offset_reg[8]  ( .D(n4404), .CLK(clk), .Q(ID_imm_offset[8]), 
        .QN(n3698) );
  DFFX1 \IF_IR_reg[7]  ( .D(n4403), .CLK(clk), .Q(N313), .QN(n3697) );
  DFFX1 \ID_imm_offset_reg[7]  ( .D(n4402), .CLK(clk), .Q(ID_imm_offset[7]), 
        .QN(n3696) );
  DFFX1 \IF_IR_reg[6]  ( .D(n4401), .CLK(clk), .Q(n5700), .QN(n3695) );
  DFFX1 \ID_imm_offset_reg[6]  ( .D(n4400), .CLK(clk), .Q(ID_imm_offset[6]), 
        .QN(n3694) );
  DFFX1 \ID_Rn_reg[0]  ( .D(n4399), .CLK(clk), .Q(ID_Rn[0]), .QN(n3693) );
  DFFX1 \ID_Rn_reg[1]  ( .D(n4398), .CLK(clk), .Q(ID_Rn[1]), .QN(n3692) );
  DFFX1 \ID_Rn_reg[2]  ( .D(n4397), .CLK(clk), .Q(ID_Rn[2]), .QN(n3691) );
  DFFX1 \ID_Rn_reg[3]  ( .D(n4396), .CLK(clk), .Q(ID_Rn[3]), .QN(n3690) );
  DFFX1 \ID_Rn_reg[4]  ( .D(n4395), .CLK(clk), .Q(ID_Rn[4]), .QN(n3689) );
  DFFX1 \ID_Rn_reg[5]  ( .D(n4394), .CLK(clk), .Q(ID_Rn[5]), .QN(n3688) );
  DFFX1 \ID_Rn_reg[6]  ( .D(n4393), .CLK(clk), .Q(ID_Rn[6]), .QN(n3687) );
  DFFX1 \ID_Rn_reg[7]  ( .D(n4392), .CLK(clk), .Q(ID_Rn[7]), .QN(n3686) );
  DFFX1 \ID_Rn_reg[8]  ( .D(n4391), .CLK(clk), .Q(ID_Rn[8]), .QN(n3685) );
  DFFX1 \ID_Rn_reg[9]  ( .D(n4390), .CLK(clk), .Q(ID_Rn[9]), .QN(n3684) );
  DFFX1 \ID_Rn_reg[10]  ( .D(n4389), .CLK(clk), .Q(ID_Rn[10]), .QN(n3683) );
  DFFX1 \ID_Rn_reg[11]  ( .D(n4388), .CLK(clk), .Q(ID_Rn[11]), .QN(n3682) );
  DFFX1 \ID_Rn_reg[12]  ( .D(n4387), .CLK(clk), .Q(ID_Rn[12]), .QN(n3681) );
  DFFX1 \ID_Rn_reg[13]  ( .D(n4386), .CLK(clk), .Q(ID_Rn[13]), .QN(n3680) );
  DFFX1 \ID_Rn_reg[14]  ( .D(n4385), .CLK(clk), .Q(ID_Rn[14]), .QN(n3679) );
  DFFX1 \ID_Rn_reg[15]  ( .D(n4384), .CLK(clk), .Q(ID_Rn[15]), .QN(n3678) );
  DFFX1 \ID_Rn_reg[16]  ( .D(n4383), .CLK(clk), .Q(ID_Rn[16]), .QN(n3677) );
  DFFX1 \ID_Rn_reg[17]  ( .D(n4382), .CLK(clk), .Q(ID_Rn[17]), .QN(n3676) );
  DFFX1 \ID_Rn_reg[18]  ( .D(n4381), .CLK(clk), .Q(ID_Rn[18]), .QN(n3675) );
  DFFX1 \ID_Rn_reg[19]  ( .D(n4380), .CLK(clk), .Q(ID_Rn[19]), .QN(n3674) );
  DFFX1 \ID_Rn_reg[20]  ( .D(n4379), .CLK(clk), .Q(ID_Rn[20]), .QN(n3673) );
  DFFX1 \ID_Rn_reg[21]  ( .D(n4378), .CLK(clk), .Q(ID_Rn[21]), .QN(n3672) );
  DFFX1 \ID_Rn_reg[22]  ( .D(n4377), .CLK(clk), .Q(ID_Rn[22]), .QN(n3671) );
  DFFX1 \ID_Rn_reg[23]  ( .D(n4376), .CLK(clk), .Q(ID_Rn[23]), .QN(n3670) );
  DFFX1 \ID_Rn_reg[24]  ( .D(n4375), .CLK(clk), .Q(ID_Rn[24]), .QN(n3669) );
  DFFX1 \ID_Rn_reg[25]  ( .D(n4374), .CLK(clk), .Q(ID_Rn[25]), .QN(n3668) );
  DFFX1 \ID_Rn_reg[26]  ( .D(n4373), .CLK(clk), .Q(ID_Rn[26]), .QN(n3667) );
  DFFX1 \ID_Rn_reg[27]  ( .D(n4372), .CLK(clk), .Q(ID_Rn[27]), .QN(n3666) );
  DFFX1 \ID_Rn_reg[28]  ( .D(n4371), .CLK(clk), .Q(ID_Rn[28]), .QN(n3665) );
  DFFX1 \ID_Rn_reg[29]  ( .D(n4370), .CLK(clk), .Q(ID_Rn[29]), .QN(n3664) );
  DFFX1 \ID_Rn_reg[30]  ( .D(n4369), .CLK(clk), .Q(ID_Rn[30]), .QN(n3663) );
  DFFX1 \ID_Rn_reg[31]  ( .D(n4368), .CLK(clk), .Q(ID_Rn[31]), .QN(n3662) );
  DFFX1 \ID_Rd_reg[31]  ( .D(n4367), .CLK(clk), .Q(N4141), .QN(n3661) );
  DFFX1 \ID_Rd_reg[30]  ( .D(n4366), .CLK(clk), .Q(ID_Rd[30]), .QN(n3660) );
  DFFX1 \ID_Rd_reg[29]  ( .D(n4365), .CLK(clk), .Q(ID_Rd[29]), .QN(n3659) );
  DFFX1 \ID_Rd_reg[28]  ( .D(n4364), .CLK(clk), .Q(ID_Rd[28]), .QN(n3658) );
  DFFX1 \ID_Rd_reg[27]  ( .D(n4363), .CLK(clk), .Q(ID_Rd[27]), .QN(n3657) );
  DFFX1 \ID_Rd_reg[26]  ( .D(n4362), .CLK(clk), .Q(ID_Rd[26]), .QN(n3656) );
  DFFX1 \ID_Rd_reg[25]  ( .D(n4361), .CLK(clk), .Q(ID_Rd[25]), .QN(n3655) );
  DFFX1 \ID_Rd_reg[24]  ( .D(n4360), .CLK(clk), .Q(ID_Rd[24]), .QN(n3654) );
  DFFX1 \ID_Rd_reg[23]  ( .D(n4359), .CLK(clk), .Q(ID_Rd[23]), .QN(n3653) );
  DFFX1 \ID_Rd_reg[22]  ( .D(n4358), .CLK(clk), .Q(ID_Rd[22]), .QN(n3652) );
  DFFX1 \ID_Rd_reg[21]  ( .D(n4357), .CLK(clk), .Q(ID_Rd[21]), .QN(n3651) );
  DFFX1 \ID_Rd_reg[20]  ( .D(n4356), .CLK(clk), .Q(ID_Rd[20]), .QN(n3650) );
  DFFX1 \ID_Rd_reg[19]  ( .D(n4355), .CLK(clk), .Q(ID_Rd[19]), .QN(n3649) );
  DFFX1 \ID_Rd_reg[18]  ( .D(n4354), .CLK(clk), .Q(ID_Rd[18]), .QN(n3648) );
  DFFX1 \ID_Rd_reg[17]  ( .D(n4353), .CLK(clk), .Q(ID_Rd[17]), .QN(n3647) );
  DFFX1 \ID_Rd_reg[16]  ( .D(n4352), .CLK(clk), .Q(ID_Rd[16]), .QN(n3646) );
  DFFX1 \ID_Rd_reg[15]  ( .D(n4351), .CLK(clk), .Q(ID_Rd[15]), .QN(n3645) );
  DFFX1 \ID_Rd_reg[14]  ( .D(n4350), .CLK(clk), .Q(ID_Rd[14]), .QN(n3644) );
  DFFX1 \ID_Rd_reg[13]  ( .D(n4349), .CLK(clk), .Q(ID_Rd[13]), .QN(n3643) );
  DFFX1 \ID_Rd_reg[12]  ( .D(n4348), .CLK(clk), .Q(ID_Rd[12]), .QN(n3642) );
  DFFX1 \ID_Rd_reg[11]  ( .D(n4347), .CLK(clk), .Q(ID_Rd[11]), .QN(n3641) );
  DFFX1 \ID_Rd_reg[10]  ( .D(n4346), .CLK(clk), .Q(ID_Rd[10]), .QN(n3640) );
  DFFX1 \ID_Rd_reg[9]  ( .D(n4345), .CLK(clk), .Q(ID_Rd[9]), .QN(n3639) );
  DFFX1 \ID_Rd_reg[8]  ( .D(n4344), .CLK(clk), .Q(ID_Rd[8]), .QN(n3638) );
  DFFX1 \ID_Rd_reg[7]  ( .D(n4343), .CLK(clk), .Q(ID_Rd[7]), .QN(n3637) );
  DFFX1 \ID_Rd_reg[6]  ( .D(n4342), .CLK(clk), .Q(ID_Rd[6]), .QN(n3636) );
  DFFX1 \ID_Rd_reg[5]  ( .D(n4341), .CLK(clk), .Q(ID_Rd[5]), .QN(n3635) );
  DFFX1 \ID_Rd_reg[4]  ( .D(n4340), .CLK(clk), .Q(ID_Rd[4]), .QN(n3634) );
  DFFX1 \ID_Rd_reg[3]  ( .D(n4339), .CLK(clk), .Q(ID_Rd[3]), .QN(n3633) );
  DFFX1 \ID_Rd_reg[2]  ( .D(n4338), .CLK(clk), .Q(ID_Rd[2]), .QN(n3632) );
  DFFX1 \ID_Rd_reg[1]  ( .D(n4337), .CLK(clk), .Q(ID_Rd[1]), .QN(n3631) );
  DFFX1 \ID_Rd_reg[0]  ( .D(n4336), .CLK(clk), .Q(ID_Rd[0]), .QN(n3630) );
  DFFX1 \ID_Rm_Rs_reg[4]  ( .D(n4331), .CLK(clk), .Q(ID_Rm_Rs[4]), .QN(n4481)
         );
  DFFX1 \ID_Rm_Rs_reg[5]  ( .D(n4330), .CLK(clk), .Q(ID_Rm_Rs[5]), .QN(n4480)
         );
  DFFX1 \ID_Rm_Rs_reg[6]  ( .D(n4329), .CLK(clk), .Q(ID_Rm_Rs[6]), .QN(n4479)
         );
  DFFX1 \ID_Rm_Rs_reg[7]  ( .D(n4328), .CLK(clk), .Q(ID_Rm_Rs[7]), .QN(n4478)
         );
  DFFX1 \ID_Rm_Rs_reg[8]  ( .D(n4327), .CLK(clk), .Q(ID_Rm_Rs[8]), .QN(n4477)
         );
  DFFX1 \ID_Rm_Rs_reg[9]  ( .D(n4326), .CLK(clk), .Q(ID_Rm_Rs[9]), .QN(n4476)
         );
  DFFX1 \ID_Rm_Rs_reg[10]  ( .D(n4325), .CLK(clk), .Q(ID_Rm_Rs[10]), .QN(n4475) );
  DFFX1 \ID_Rm_Rs_reg[11]  ( .D(n4324), .CLK(clk), .Q(ID_Rm_Rs[11]), .QN(n4474) );
  DFFX1 \ID_Rm_Rs_reg[12]  ( .D(n4323), .CLK(clk), .Q(ID_Rm_Rs[12]), .QN(n4473) );
  DFFX1 \ID_Rm_Rs_reg[13]  ( .D(n4322), .CLK(clk), .Q(ID_Rm_Rs[13]), .QN(n4472) );
  DFFX1 \ID_Rm_Rs_reg[14]  ( .D(n4321), .CLK(clk), .Q(ID_Rm_Rs[14]), .QN(n4471) );
  DFFX1 \ID_Rm_Rs_reg[15]  ( .D(n4320), .CLK(clk), .Q(ID_Rm_Rs[15]), .QN(n4470) );
  DFFX1 \ID_Rm_Rs_reg[16]  ( .D(n4319), .CLK(clk), .Q(ID_Rm_Rs[16]), .QN(n4469) );
  DFFX1 \ID_Rm_Rs_reg[17]  ( .D(n4318), .CLK(clk), .Q(ID_Rm_Rs[17]), .QN(n4468) );
  DFFX1 \ID_Rm_Rs_reg[18]  ( .D(n4317), .CLK(clk), .Q(ID_Rm_Rs[18]), .QN(n4467) );
  DFFX1 \ID_Rm_Rs_reg[19]  ( .D(n4316), .CLK(clk), .Q(ID_Rm_Rs[19]), .QN(n4466) );
  DFFX1 \ID_Rm_Rs_reg[20]  ( .D(n4315), .CLK(clk), .Q(ID_Rm_Rs[20]), .QN(n4465) );
  DFFX1 \ID_Rm_Rs_reg[21]  ( .D(n4314), .CLK(clk), .Q(ID_Rm_Rs[21]), .QN(n4464) );
  DFFX1 \ID_Rm_Rs_reg[22]  ( .D(n4313), .CLK(clk), .Q(ID_Rm_Rs[22]), .QN(n4463) );
  DFFX1 \ID_Rm_Rs_reg[23]  ( .D(n4312), .CLK(clk), .Q(ID_Rm_Rs[23]), .QN(n4462) );
  DFFX1 \ID_Rm_Rs_reg[24]  ( .D(n4311), .CLK(clk), .Q(ID_Rm_Rs[24]), .QN(n4461) );
  DFFX1 \ID_Rm_Rs_reg[25]  ( .D(n4310), .CLK(clk), .Q(ID_Rm_Rs[25]), .QN(n4460) );
  DFFX1 \ID_Rm_Rs_reg[26]  ( .D(n4309), .CLK(clk), .Q(ID_Rm_Rs[26]), .QN(n4459) );
  DFFX1 \ID_Rm_Rs_reg[27]  ( .D(n4308), .CLK(clk), .Q(ID_Rm_Rs[27]), .QN(n4458) );
  DFFX1 \ID_Rm_Rs_reg[28]  ( .D(n4307), .CLK(clk), .Q(ID_Rm_Rs[28]), .QN(n4457) );
  DFFX1 \ID_Rm_Rs_reg[29]  ( .D(n4306), .CLK(clk), .Q(ID_Rm_Rs[29]), .QN(n4456) );
  DFFX1 \ID_Rm_Rs_reg[30]  ( .D(n4305), .CLK(clk), .Q(ID_Rm_Rs[30]), .QN(n4455) );
  DFFX1 \ID_Rm_Rs_reg[31]  ( .D(n4304), .CLK(clk), .Q(N3016), .QN(n4454) );
  DFFX1 \IF_IR_reg[5]  ( .D(n4303), .CLK(clk), .Q(N308), .QN(n9195) );
  DFFX1 \ID_imm_offset_reg[5]  ( .D(n4302), .CLK(clk), .Q(ID_imm_offset[5]), 
        .QN(n3629) );
  DFFX1 \IF_IR_reg[4]  ( .D(n4301), .CLK(clk), .Q(N307), .QN(n9196) );
  DFFX1 \ID_imm_offset_reg[4]  ( .D(n4300), .CLK(clk), .Q(ID_imm_offset[4]), 
        .QN(n3628) );
  DFFX1 \IF_IR_reg[3]  ( .D(n4299), .CLK(clk), .Q(n5699), .QN(n9197) );
  DFFX1 \IF_IR_reg[2]  ( .D(n4297), .CLK(clk), .Q(N311), .QN(n9192) );
  DFFX1 \ID_Rd_code_reg[2]  ( .D(n4295), .CLK(clk), .Q(n9165) );
  DFFX1 \IF_IR_reg[1]  ( .D(n4294), .CLK(clk), .Q(N310), .QN(n9193) );
  DFFX1 \ID_Rd_code_reg[1]  ( .D(n4292), .CLK(clk), .Q(n9164) );
  DFFX1 \IF_IR_reg[0]  ( .D(n4291), .CLK(clk), .Q(n5698), .QN(n9194) );
  DFFX1 \ID_Rd_code_reg[0]  ( .D(n4289), .CLK(clk), .Q(n9163) );
  DFFX1 \EX_opcode_reg[4]  ( .D(n4288), .CLK(clk), .Q(n9181), .QN(n5703) );
  DFFX1 \EX_opcode_reg[2]  ( .D(n4287), .CLK(clk), .Q(n9183), .QN(n5693) );
  DFFX1 \EX_opcode_reg[1]  ( .D(n4286), .CLK(clk), .Q(n9179), .QN(n5688) );
  DFFX1 \EX_opcode_reg[0]  ( .D(n4285), .CLK(clk), .Q(n9180), .QN(n5708) );
  DFFX1 \EX_opcode_reg[3]  ( .D(n4284), .CLK(clk), .Q(n9184), .QN(n5710) );
  DFFX1 \EX_opcode_reg[5]  ( .D(n4283), .CLK(clk), .Q(n9182), .QN(n5707) );
  DFFX1 \EX_Rd_code_reg[0]  ( .D(n4282), .CLK(clk), .Q(n9162), .QN(n5704) );
  DFFX1 \EX_Rd_code_reg[1]  ( .D(n4281), .CLK(clk), .Q(n9161), .QN(n5691) );
  DFFX1 \EX_Rd_code_reg[2]  ( .D(n4280), .CLK(clk), .Q(n9160) );
  DFFX1 \DR_reg[0]  ( .D(n4279), .CLK(clk), .Q(n9199) );
  DFFX1 \DR_reg[1]  ( .D(n4278), .CLK(clk), .Q(n9200) );
  DFFX1 \DR_reg[2]  ( .D(n4277), .CLK(clk), .Q(n9201) );
  DFFX1 \DR_reg[3]  ( .D(n4276), .CLK(clk), .Q(n9202) );
  DFFX1 \DR_reg[4]  ( .D(n4275), .CLK(clk), .Q(n9203) );
  DFFX1 \DR_reg[5]  ( .D(n4274), .CLK(clk), .Q(n9204) );
  DFFX1 \DR_reg[6]  ( .D(n4273), .CLK(clk), .Q(n9205) );
  DFFX1 \DR_reg[7]  ( .D(n4272), .CLK(clk), .Q(n9206) );
  DFFX1 \DR_reg[8]  ( .D(n4271), .CLK(clk), .Q(n9207) );
  DFFX1 \DR_reg[9]  ( .D(n4270), .CLK(clk), .Q(n9208) );
  DFFX1 \DR_reg[10]  ( .D(n4269), .CLK(clk), .Q(n9209) );
  DFFX1 \DR_reg[11]  ( .D(n4268), .CLK(clk), .Q(n9210) );
  DFFX1 \DR_reg[12]  ( .D(n4267), .CLK(clk), .Q(n9211) );
  DFFX1 \DR_reg[13]  ( .D(n4266), .CLK(clk), .Q(n9212) );
  DFFX1 \DR_reg[14]  ( .D(n4265), .CLK(clk), .Q(n9213) );
  DFFX1 \DR_reg[15]  ( .D(n4264), .CLK(clk), .Q(n9214) );
  DFFX1 \DR_reg[16]  ( .D(n4263), .CLK(clk), .Q(n9215) );
  DFFX1 \DR_reg[17]  ( .D(n4262), .CLK(clk), .Q(n9216) );
  DFFX1 \DR_reg[18]  ( .D(n4261), .CLK(clk), .Q(n9217) );
  DFFX1 \DR_reg[19]  ( .D(n4260), .CLK(clk), .Q(n9218) );
  DFFX1 \DR_reg[20]  ( .D(n4259), .CLK(clk), .Q(n9219) );
  DFFX1 \DR_reg[21]  ( .D(n4258), .CLK(clk), .Q(n9220) );
  DFFX1 \DR_reg[22]  ( .D(n4257), .CLK(clk), .Q(n9221) );
  DFFX1 \DR_reg[23]  ( .D(n4256), .CLK(clk), .Q(n9222) );
  DFFX1 \DR_reg[24]  ( .D(n4255), .CLK(clk), .Q(n9223) );
  DFFX1 \DR_reg[25]  ( .D(n4254), .CLK(clk), .Q(n9224) );
  DFFX1 \DR_reg[26]  ( .D(n4253), .CLK(clk), .Q(n9225) );
  DFFX1 \DR_reg[27]  ( .D(n4252), .CLK(clk), .Q(n9226) );
  DFFX1 \DR_reg[28]  ( .D(n4251), .CLK(clk), .Q(n9227) );
  DFFX1 \DR_reg[29]  ( .D(n4250), .CLK(clk), .Q(n9228) );
  DFFX1 \DR_reg[30]  ( .D(n4249), .CLK(clk), .Q(n9229) );
  DFFX1 \DR_reg[31]  ( .D(n4248), .CLK(clk), .Q(n9230) );
  DFFX1 \EX_imm_offset_reg[7]  ( .D(n4247), .CLK(clk), .Q(n9174), .QN(n5687)
         );
  DFFX1 \EX_imm_offset_reg[6]  ( .D(n4246), .CLK(clk), .Q(n9159), .QN(n5713)
         );
  DFFX1 \EX_imm_offset_reg[5]  ( .D(n4245), .CLK(clk), .Q(n9175), .QN(n5690)
         );
  DFFX1 \EX_imm_offset_reg[4]  ( .D(n4244), .CLK(clk), .Q(n9158), .QN(n5694)
         );
  DFFX1 \EX_imm_offset_reg[3]  ( .D(n4243), .CLK(clk), .Q(n9178) );
  DFFX1 \EX_imm_offset_reg[2]  ( .D(n4242), .CLK(clk), .Q(n9177), .QN(n5714)
         );
  DFFX1 \EX_imm_offset_reg[1]  ( .D(n4241), .CLK(clk), .Q(n9176) );
  DFFX1 \SP_reg[31]  ( .D(n4240), .CLK(clk), .Q(SP[31]) );
  DFFX1 \SP_reg[0]  ( .D(n4239), .CLK(clk), .Q(SP[0]), .QN(n3574) );
  DFFX1 \SP_reg[1]  ( .D(n4238), .CLK(clk), .Q(SP[1]), .QN(n3573) );
  DFFX1 \SP_reg[2]  ( .D(n4237), .CLK(clk), .Q(SP[2]) );
  DFFX1 \SP_reg[3]  ( .D(n4236), .CLK(clk), .Q(SP[3]) );
  DFFX1 \SP_reg[4]  ( .D(n4235), .CLK(clk), .Q(SP[4]) );
  DFFX1 \SP_reg[5]  ( .D(n4234), .CLK(clk), .Q(SP[5]) );
  DFFX1 \SP_reg[6]  ( .D(n4233), .CLK(clk), .Q(SP[6]) );
  DFFX1 \SP_reg[7]  ( .D(n4232), .CLK(clk), .Q(SP[7]) );
  DFFX1 \SP_reg[8]  ( .D(n4231), .CLK(clk), .Q(SP[8]) );
  DFFX1 \SP_reg[9]  ( .D(n4230), .CLK(clk), .Q(SP[9]) );
  DFFX1 \SP_reg[10]  ( .D(n4229), .CLK(clk), .Q(SP[10]) );
  DFFX1 \SP_reg[11]  ( .D(n4228), .CLK(clk), .Q(SP[11]) );
  DFFX1 \SP_reg[12]  ( .D(n4227), .CLK(clk), .Q(SP[12]) );
  DFFX1 \SP_reg[13]  ( .D(n4226), .CLK(clk), .Q(SP[13]) );
  DFFX1 \SP_reg[14]  ( .D(n4225), .CLK(clk), .Q(SP[14]) );
  DFFX1 \SP_reg[15]  ( .D(n4224), .CLK(clk), .Q(SP[15]) );
  DFFX1 \SP_reg[16]  ( .D(n4223), .CLK(clk), .Q(SP[16]) );
  DFFX1 \SP_reg[17]  ( .D(n4222), .CLK(clk), .Q(SP[17]) );
  DFFX1 \SP_reg[18]  ( .D(n4221), .CLK(clk), .Q(SP[18]) );
  DFFX1 \SP_reg[19]  ( .D(n4220), .CLK(clk), .Q(SP[19]) );
  DFFX1 \SP_reg[20]  ( .D(n4219), .CLK(clk), .Q(SP[20]) );
  DFFX1 \SP_reg[21]  ( .D(n4218), .CLK(clk), .Q(SP[21]) );
  DFFX1 \SP_reg[22]  ( .D(n4217), .CLK(clk), .Q(SP[22]) );
  DFFX1 \SP_reg[23]  ( .D(n4216), .CLK(clk), .Q(SP[23]) );
  DFFX1 \SP_reg[24]  ( .D(n4215), .CLK(clk), .Q(SP[24]) );
  DFFX1 \SP_reg[25]  ( .D(n4214), .CLK(clk), .Q(SP[25]) );
  DFFX1 \SP_reg[26]  ( .D(n4213), .CLK(clk), .Q(SP[26]) );
  DFFX1 \SP_reg[27]  ( .D(n4212), .CLK(clk), .Q(SP[27]) );
  DFFX1 \SP_reg[28]  ( .D(n4211), .CLK(clk), .Q(SP[28]) );
  DFFX1 \SP_reg[29]  ( .D(n4210), .CLK(clk), .Q(SP[29]) );
  DFFX1 \SP_reg[30]  ( .D(n4209), .CLK(clk), .Q(SP[30]) );
  DFFX1 \ALU_out_reg[32]  ( .D(n4208), .CLK(clk), .Q(n9157) );
  DFFX1 \ALU_out_reg[0]  ( .D(n4207), .CLK(clk), .Q(n9156) );
  DFFX1 \data_address_reg[0]  ( .D(n4206), .CLK(clk), .Q(data_address[0]) );
  DFFX1 \ALU_out_reg[1]  ( .D(n4205), .CLK(clk), .Q(n9155) );
  DFFX1 \data_address_reg[1]  ( .D(n4204), .CLK(clk), .Q(data_address[1]) );
  DFFX1 \ALU_out_reg[2]  ( .D(n4203), .CLK(clk), .Q(n9154) );
  DFFX1 \data_address_reg[2]  ( .D(n4202), .CLK(clk), .Q(data_address[2]) );
  DFFX1 \ALU_out_reg[3]  ( .D(n4201), .CLK(clk), .Q(n9153) );
  DFFX1 \data_address_reg[3]  ( .D(n4200), .CLK(clk), .Q(data_address[3]) );
  DFFX1 \ALU_out_reg[4]  ( .D(n4199), .CLK(clk), .Q(n9152) );
  DFFX1 \data_address_reg[4]  ( .D(n4198), .CLK(clk), .Q(data_address[4]) );
  DFFX1 \ALU_out_reg[5]  ( .D(n4197), .CLK(clk), .Q(n9151) );
  DFFX1 \data_address_reg[5]  ( .D(n4196), .CLK(clk), .Q(data_address[5]) );
  DFFX1 \ALU_out_reg[6]  ( .D(n4195), .CLK(clk), .Q(n9150) );
  DFFX1 \data_address_reg[6]  ( .D(n4194), .CLK(clk), .Q(data_address[6]) );
  DFFX1 \ALU_out_reg[7]  ( .D(n4193), .CLK(clk), .Q(n9149) );
  DFFX1 \data_address_reg[7]  ( .D(n4192), .CLK(clk), .Q(data_address[7]) );
  DFFX1 \ALU_out_reg[8]  ( .D(n4191), .CLK(clk), .Q(n9148) );
  DFFX1 \data_address_reg[8]  ( .D(n4190), .CLK(clk), .Q(data_address[8]) );
  DFFX1 \ALU_out_reg[9]  ( .D(n4189), .CLK(clk), .Q(n9147) );
  DFFX1 \data_address_reg[9]  ( .D(n4188), .CLK(clk), .Q(data_address[9]) );
  DFFX1 \ALU_out_reg[10]  ( .D(n4187), .CLK(clk), .Q(n9146) );
  DFFX1 \data_address_reg[10]  ( .D(n4186), .CLK(clk), .Q(data_address[10]) );
  DFFX1 \ALU_out_reg[11]  ( .D(n4185), .CLK(clk), .Q(n9145) );
  DFFX1 \data_address_reg[11]  ( .D(n4184), .CLK(clk), .Q(data_address[11]) );
  DFFX1 \ALU_out_reg[12]  ( .D(n4183), .CLK(clk), .Q(n9144) );
  DFFX1 \data_address_reg[12]  ( .D(n4182), .CLK(clk), .Q(data_address[12]) );
  DFFX1 \ALU_out_reg[13]  ( .D(n4181), .CLK(clk), .Q(n9143) );
  DFFX1 \data_address_reg[13]  ( .D(n4180), .CLK(clk), .Q(data_address[13]) );
  DFFX1 \ALU_out_reg[14]  ( .D(n4179), .CLK(clk), .Q(n9142) );
  DFFX1 \data_address_reg[14]  ( .D(n4178), .CLK(clk), .Q(data_address[14]) );
  DFFX1 \ALU_out_reg[15]  ( .D(n4177), .CLK(clk), .Q(n9141) );
  DFFX1 \data_address_reg[15]  ( .D(n4176), .CLK(clk), .Q(data_address[15]) );
  DFFX1 \ALU_out_reg[16]  ( .D(n4175), .CLK(clk), .Q(n9140) );
  DFFX1 \data_address_reg[16]  ( .D(n4174), .CLK(clk), .Q(data_address[16]) );
  DFFX1 \ALU_out_reg[17]  ( .D(n4173), .CLK(clk), .Q(n9139) );
  DFFX1 \data_address_reg[17]  ( .D(n4172), .CLK(clk), .Q(data_address[17]) );
  DFFX1 \ALU_out_reg[18]  ( .D(n4171), .CLK(clk), .Q(n9138) );
  DFFX1 \data_address_reg[18]  ( .D(n4170), .CLK(clk), .Q(data_address[18]) );
  DFFX1 \ALU_out_reg[19]  ( .D(n4169), .CLK(clk), .Q(n9137) );
  DFFX1 \data_address_reg[19]  ( .D(n4168), .CLK(clk), .Q(data_address[19]) );
  DFFX1 \ALU_out_reg[20]  ( .D(n4167), .CLK(clk), .Q(n9136) );
  DFFX1 \data_address_reg[20]  ( .D(n4166), .CLK(clk), .Q(data_address[20]) );
  DFFX1 \ALU_out_reg[21]  ( .D(n4165), .CLK(clk), .Q(n9135) );
  DFFX1 \data_address_reg[21]  ( .D(n4164), .CLK(clk), .Q(data_address[21]) );
  DFFX1 \ALU_out_reg[22]  ( .D(n4163), .CLK(clk), .Q(n9134) );
  DFFX1 \data_address_reg[22]  ( .D(n4162), .CLK(clk), .Q(data_address[22]) );
  DFFX1 \ALU_out_reg[23]  ( .D(n4161), .CLK(clk), .Q(n9133) );
  DFFX1 \data_address_reg[23]  ( .D(n4160), .CLK(clk), .Q(data_address[23]) );
  DFFX1 \ALU_out_reg[24]  ( .D(n4159), .CLK(clk), .Q(n9132) );
  DFFX1 \data_address_reg[24]  ( .D(n4158), .CLK(clk), .Q(data_address[24]) );
  DFFX1 \ALU_out_reg[25]  ( .D(n4157), .CLK(clk), .Q(n9131) );
  DFFX1 \data_address_reg[25]  ( .D(n4156), .CLK(clk), .Q(data_address[25]) );
  DFFX1 \ALU_out_reg[26]  ( .D(n4155), .CLK(clk), .Q(n9130) );
  DFFX1 \data_address_reg[26]  ( .D(n4154), .CLK(clk), .Q(data_address[26]) );
  DFFX1 \ALU_out_reg[27]  ( .D(n4153), .CLK(clk), .Q(n9129) );
  DFFX1 \data_address_reg[27]  ( .D(n4152), .CLK(clk), .Q(data_address[27]) );
  DFFX1 \ALU_out_reg[28]  ( .D(n4151), .CLK(clk), .Q(n9128) );
  DFFX1 \data_address_reg[28]  ( .D(n4150), .CLK(clk), .Q(data_address[28]) );
  DFFX1 \ALU_out_reg[29]  ( .D(n4149), .CLK(clk), .Q(n9127) );
  DFFX1 \data_address_reg[29]  ( .D(n4148), .CLK(clk), .Q(data_address[29]) );
  DFFX1 \ALU_out_reg[30]  ( .D(n4147), .CLK(clk), .Q(n9126) );
  DFFX1 \data_address_reg[30]  ( .D(n4146), .CLK(clk), .Q(data_address[30]) );
  DFFX1 \ALU_out_reg[31]  ( .D(n4145), .CLK(clk), .Q(n9125) );
  DFFX1 \data_address_reg[31]  ( .D(n4144), .CLK(clk), .Q(data_address[31]) );
  DFFX1 N_Flag_reg ( .D(n4143), .CLK(clk), .Q(n9124) );
  DFFX1 Z_Flag_reg ( .D(n4142), .CLK(clk), .Q(n9123) );
  DFFX1 C_Flag_reg ( .D(n4141), .CLK(clk), .Q(n9173), .QN(n4486) );
  DFFX1 \branch_target_reg[0]  ( .D(n4140), .CLK(clk), .Q(n9122) );
  DFFX1 \branch_target_reg[1]  ( .D(n4139), .CLK(clk), .Q(n9121) );
  DFFX1 \LR_reg[1]  ( .D(n4138), .CLK(clk), .Q(n9120) );
  DFFX1 \branch_target_reg[2]  ( .D(n4137), .CLK(clk), .Q(n9119) );
  DFFX1 \LR_reg[2]  ( .D(n4136), .CLK(clk), .Q(n9118) );
  DFFX1 \branch_target_reg[3]  ( .D(n4135), .CLK(clk), .Q(n9117) );
  DFFX1 \LR_reg[3]  ( .D(n4134), .CLK(clk), .Q(n9116) );
  DFFX1 \branch_target_reg[4]  ( .D(n4133), .CLK(clk), .Q(n9115) );
  DFFX1 \LR_reg[4]  ( .D(n4132), .CLK(clk), .Q(n9114) );
  DFFX1 \branch_target_reg[5]  ( .D(n4131), .CLK(clk), .Q(n9113) );
  DFFX1 \LR_reg[5]  ( .D(n4130), .CLK(clk), .Q(n9112) );
  DFFX1 \branch_target_reg[6]  ( .D(n4129), .CLK(clk), .Q(n9111) );
  DFFX1 \LR_reg[6]  ( .D(n4128), .CLK(clk), .Q(n9110) );
  DFFX1 \branch_target_reg[7]  ( .D(n4127), .CLK(clk), .Q(n9109) );
  DFFX1 \LR_reg[7]  ( .D(n4126), .CLK(clk), .Q(n9108) );
  DFFX1 \branch_target_reg[8]  ( .D(n4125), .CLK(clk), .Q(n9107) );
  DFFX1 \LR_reg[8]  ( .D(n4124), .CLK(clk), .Q(n9106) );
  DFFX1 \branch_target_reg[9]  ( .D(n4123), .CLK(clk), .Q(n9105) );
  DFFX1 \LR_reg[9]  ( .D(n4122), .CLK(clk), .Q(n9104) );
  DFFX1 \branch_target_reg[10]  ( .D(n4121), .CLK(clk), .Q(n9103) );
  DFFX1 \LR_reg[10]  ( .D(n4120), .CLK(clk), .Q(n9102) );
  DFFX1 \branch_target_reg[11]  ( .D(n4119), .CLK(clk), .Q(n9101) );
  DFFX1 \LR_reg[11]  ( .D(n4118), .CLK(clk), .Q(n9100) );
  DFFX1 \branch_target_reg[12]  ( .D(n4117), .CLK(clk), .Q(n9099) );
  DFFX1 \LR_reg[12]  ( .D(n4116), .CLK(clk), .Q(n9098) );
  DFFX1 \branch_target_reg[13]  ( .D(n4115), .CLK(clk), .Q(n9097) );
  DFFX1 \LR_reg[13]  ( .D(n4114), .CLK(clk), .Q(n9096) );
  DFFX1 \branch_target_reg[14]  ( .D(n4113), .CLK(clk), .Q(n9095) );
  DFFX1 \LR_reg[14]  ( .D(n4112), .CLK(clk), .Q(n9094) );
  DFFX1 \branch_target_reg[15]  ( .D(n4111), .CLK(clk), .Q(n9093) );
  DFFX1 \LR_reg[15]  ( .D(n4110), .CLK(clk), .Q(n9092) );
  DFFX1 \branch_target_reg[16]  ( .D(n4109), .CLK(clk), .Q(n9091) );
  DFFX1 \LR_reg[16]  ( .D(n4108), .CLK(clk), .Q(n9090) );
  DFFX1 \branch_target_reg[17]  ( .D(n4107), .CLK(clk), .Q(n9089) );
  DFFX1 \LR_reg[17]  ( .D(n4106), .CLK(clk), .Q(n9088) );
  DFFX1 \branch_target_reg[18]  ( .D(n4105), .CLK(clk), .Q(n9087) );
  DFFX1 \LR_reg[18]  ( .D(n4104), .CLK(clk), .Q(n9086) );
  DFFX1 \branch_target_reg[19]  ( .D(n4103), .CLK(clk), .Q(n9085) );
  DFFX1 \LR_reg[19]  ( .D(n4102), .CLK(clk), .Q(n9084) );
  DFFX1 \branch_target_reg[20]  ( .D(n4101), .CLK(clk), .Q(n9083) );
  DFFX1 \LR_reg[20]  ( .D(n4100), .CLK(clk), .Q(n9082) );
  DFFX1 \branch_target_reg[21]  ( .D(n4099), .CLK(clk), .Q(n9081) );
  DFFX1 \LR_reg[21]  ( .D(n4098), .CLK(clk), .Q(n9080) );
  DFFX1 \branch_target_reg[22]  ( .D(n4097), .CLK(clk), .Q(n9079) );
  DFFX1 \LR_reg[22]  ( .D(n4096), .CLK(clk), .Q(n9078) );
  DFFX1 \branch_target_reg[23]  ( .D(n4095), .CLK(clk), .Q(n9077) );
  DFFX1 \LR_reg[23]  ( .D(n4094), .CLK(clk), .Q(n9076) );
  DFFX1 \branch_target_reg[24]  ( .D(n4093), .CLK(clk), .Q(n9075) );
  DFFX1 \LR_reg[24]  ( .D(n4092), .CLK(clk), .Q(n9074) );
  DFFX1 \branch_target_reg[25]  ( .D(n4091), .CLK(clk), .Q(n9073) );
  DFFX1 \LR_reg[25]  ( .D(n4090), .CLK(clk), .Q(n9072) );
  DFFX1 \branch_target_reg[26]  ( .D(n4089), .CLK(clk), .Q(n9071) );
  DFFX1 \LR_reg[26]  ( .D(n4088), .CLK(clk), .Q(n9070) );
  DFFX1 \branch_target_reg[27]  ( .D(n4087), .CLK(clk), .Q(n9069) );
  DFFX1 \LR_reg[27]  ( .D(n4086), .CLK(clk), .Q(n9068) );
  DFFX1 \branch_target_reg[28]  ( .D(n4085), .CLK(clk), .Q(n9067) );
  DFFX1 \LR_reg[28]  ( .D(n4084), .CLK(clk), .Q(n9066) );
  DFFX1 \branch_target_reg[29]  ( .D(n4083), .CLK(clk), .Q(n9065) );
  DFFX1 \LR_reg[29]  ( .D(n4082), .CLK(clk), .Q(n9064) );
  DFFX1 \branch_target_reg[30]  ( .D(n4081), .CLK(clk), .Q(n9063) );
  DFFX1 \LR_reg[30]  ( .D(n4080), .CLK(clk), .Q(n9062) );
  DFFX1 \branch_target_reg[31]  ( .D(n4079), .CLK(clk), .Q(n9061) );
  DFFX1 \IF_PC_reg[31]  ( .D(n4078), .CLK(clk), .Q(IF_PC[31]) );
  DFFX1 \IF_PC_reg[0]  ( .D(n4077), .CLK(clk), .Q(IF_PC[0]) );
  DFFX1 \IF_PC_reg[1]  ( .D(n4076), .CLK(clk), .Q(IF_PC[1]) );
  DFFX1 \IF_PC_reg[2]  ( .D(n4075), .CLK(clk), .Q(IF_PC[2]) );
  DFFX1 \IF_PC_reg[3]  ( .D(n4074), .CLK(clk), .Q(IF_PC[3]) );
  DFFX1 \IF_PC_reg[4]  ( .D(n4073), .CLK(clk), .Q(IF_PC[4]) );
  DFFX1 \IF_PC_reg[5]  ( .D(n4072), .CLK(clk), .Q(IF_PC[5]) );
  DFFX1 \IF_PC_reg[6]  ( .D(n4071), .CLK(clk), .Q(IF_PC[6]) );
  DFFX1 \IF_PC_reg[7]  ( .D(n4070), .CLK(clk), .Q(IF_PC[7]) );
  DFFX1 \IF_PC_reg[8]  ( .D(n4069), .CLK(clk), .Q(IF_PC[8]) );
  DFFX1 \IF_PC_reg[9]  ( .D(n4068), .CLK(clk), .Q(IF_PC[9]) );
  DFFX1 \IF_PC_reg[10]  ( .D(n4067), .CLK(clk), .Q(IF_PC[10]) );
  DFFX1 \IF_PC_reg[11]  ( .D(n4066), .CLK(clk), .Q(IF_PC[11]) );
  DFFX1 \IF_PC_reg[12]  ( .D(n4065), .CLK(clk), .Q(IF_PC[12]) );
  DFFX1 \IF_PC_reg[13]  ( .D(n4064), .CLK(clk), .Q(IF_PC[13]) );
  DFFX1 \IF_PC_reg[14]  ( .D(n4063), .CLK(clk), .Q(IF_PC[14]) );
  DFFX1 \IF_PC_reg[15]  ( .D(n4062), .CLK(clk), .Q(IF_PC[15]) );
  DFFX1 \IF_PC_reg[16]  ( .D(n4061), .CLK(clk), .Q(IF_PC[16]) );
  DFFX1 \IF_PC_reg[17]  ( .D(n4060), .CLK(clk), .Q(IF_PC[17]) );
  DFFX1 \IF_PC_reg[18]  ( .D(n4059), .CLK(clk), .Q(IF_PC[18]) );
  DFFX1 \IF_PC_reg[19]  ( .D(n4058), .CLK(clk), .Q(IF_PC[19]) );
  DFFX1 \IF_PC_reg[20]  ( .D(n4057), .CLK(clk), .Q(IF_PC[20]) );
  DFFX1 \IF_PC_reg[21]  ( .D(n4056), .CLK(clk), .Q(IF_PC[21]) );
  DFFX1 \IF_PC_reg[22]  ( .D(n4055), .CLK(clk), .Q(IF_PC[22]) );
  DFFX1 \IF_PC_reg[23]  ( .D(n4054), .CLK(clk), .Q(IF_PC[23]) );
  DFFX1 \IF_PC_reg[24]  ( .D(n4053), .CLK(clk), .Q(IF_PC[24]) );
  DFFX1 \IF_PC_reg[25]  ( .D(n4052), .CLK(clk), .Q(IF_PC[25]) );
  DFFX1 \IF_PC_reg[26]  ( .D(n4051), .CLK(clk), .Q(IF_PC[26]) );
  DFFX1 \IF_PC_reg[27]  ( .D(n4050), .CLK(clk), .Q(IF_PC[27]) );
  DFFX1 \IF_PC_reg[28]  ( .D(n4049), .CLK(clk), .Q(IF_PC[28]) );
  DFFX1 \IF_PC_reg[29]  ( .D(n4048), .CLK(clk), .Q(IF_PC[29]) );
  DFFX1 \IF_PC_reg[30]  ( .D(n4047), .CLK(clk), .Q(IF_PC[30]) );
  DFFX1 \EX_ALU_out_reg[0]  ( .D(n4046), .CLK(clk), .Q(n9060) );
  DFFX1 \EX_ALU_out_reg[1]  ( .D(n4045), .CLK(clk), .Q(n9059) );
  DFFX1 \EX_ALU_out_reg[2]  ( .D(n4044), .CLK(clk), .Q(n9058) );
  DFFX1 \EX_ALU_out_reg[3]  ( .D(n4043), .CLK(clk), .Q(n9057) );
  DFFX1 \EX_ALU_out_reg[4]  ( .D(n4042), .CLK(clk), .Q(n9056) );
  DFFX1 \EX_ALU_out_reg[5]  ( .D(n4041), .CLK(clk), .Q(n9055) );
  DFFX1 \EX_ALU_out_reg[6]  ( .D(n4040), .CLK(clk), .Q(n9054) );
  DFFX1 \EX_ALU_out_reg[7]  ( .D(n4039), .CLK(clk), .Q(n9053) );
  DFFX1 \EX_ALU_out_reg[8]  ( .D(n4038), .CLK(clk), .Q(n9052) );
  DFFX1 \EX_ALU_out_reg[9]  ( .D(n4037), .CLK(clk), .Q(n9051) );
  DFFX1 \EX_ALU_out_reg[10]  ( .D(n4036), .CLK(clk), .Q(n9050) );
  DFFX1 \EX_ALU_out_reg[11]  ( .D(n4035), .CLK(clk), .Q(n9049) );
  DFFX1 \EX_ALU_out_reg[12]  ( .D(n4034), .CLK(clk), .Q(n9048) );
  DFFX1 \EX_ALU_out_reg[13]  ( .D(n4033), .CLK(clk), .Q(n9047) );
  DFFX1 \EX_ALU_out_reg[14]  ( .D(n4032), .CLK(clk), .Q(n9046) );
  DFFX1 \EX_ALU_out_reg[15]  ( .D(n4031), .CLK(clk), .Q(n9045) );
  DFFX1 \EX_ALU_out_reg[16]  ( .D(n4030), .CLK(clk), .Q(n9044) );
  DFFX1 \EX_ALU_out_reg[17]  ( .D(n4029), .CLK(clk), .Q(n9043) );
  DFFX1 \EX_ALU_out_reg[18]  ( .D(n4028), .CLK(clk), .Q(n9042) );
  DFFX1 \EX_ALU_out_reg[19]  ( .D(n4027), .CLK(clk), .Q(n9041) );
  DFFX1 \EX_ALU_out_reg[20]  ( .D(n4026), .CLK(clk), .Q(n9040) );
  DFFX1 \EX_ALU_out_reg[21]  ( .D(n4025), .CLK(clk), .Q(n9039) );
  DFFX1 \EX_ALU_out_reg[22]  ( .D(n4024), .CLK(clk), .Q(n9038) );
  DFFX1 \EX_ALU_out_reg[23]  ( .D(n4023), .CLK(clk), .Q(n9037) );
  DFFX1 \EX_ALU_out_reg[24]  ( .D(n4022), .CLK(clk), .Q(n9036) );
  DFFX1 \EX_ALU_out_reg[25]  ( .D(n4021), .CLK(clk), .Q(n9035) );
  DFFX1 \EX_ALU_out_reg[26]  ( .D(n4020), .CLK(clk), .Q(n9034) );
  DFFX1 \EX_ALU_out_reg[27]  ( .D(n4019), .CLK(clk), .Q(n9033) );
  DFFX1 \EX_ALU_out_reg[28]  ( .D(n4018), .CLK(clk), .Q(n9032) );
  DFFX1 \EX_ALU_out_reg[29]  ( .D(n4017), .CLK(clk), .Q(n9031) );
  DFFX1 \EX_ALU_out_reg[30]  ( .D(n4016), .CLK(clk), .Q(n9030) );
  DFFX1 \EX_ALU_out_reg[31]  ( .D(n4015), .CLK(clk), .Q(n9029) );
  DFFX1 \LR_reg[31]  ( .D(n4014), .CLK(clk), .Q(n9028) );
  DFFASX1 \R_reg[7][31]  ( .D(n4013), .CLK(clk), .SETB(reset_n), .Q(\R[7][31] ) );
  DFFASX1 \R_reg[7][30]  ( .D(n4012), .CLK(clk), .SETB(reset_n), .Q(\R[7][30] ) );
  DFFASX1 \R_reg[7][29]  ( .D(n4011), .CLK(clk), .SETB(reset_n), .Q(\R[7][29] ) );
  DFFASX1 \R_reg[7][28]  ( .D(n4010), .CLK(clk), .SETB(reset_n), .Q(\R[7][28] ) );
  DFFASX1 \R_reg[7][27]  ( .D(n4009), .CLK(clk), .SETB(reset_n), .Q(\R[7][27] ) );
  DFFASX1 \R_reg[7][26]  ( .D(n4008), .CLK(clk), .SETB(reset_n), .Q(\R[7][26] ) );
  DFFASX1 \R_reg[7][25]  ( .D(n4007), .CLK(clk), .SETB(reset_n), .Q(\R[7][25] ) );
  DFFASX1 \R_reg[7][24]  ( .D(n4006), .CLK(clk), .SETB(reset_n), .Q(\R[7][24] ) );
  DFFASX1 \R_reg[7][23]  ( .D(n4005), .CLK(clk), .SETB(reset_n), .Q(\R[7][23] ) );
  DFFASX1 \R_reg[7][22]  ( .D(n4004), .CLK(clk), .SETB(reset_n), .Q(\R[7][22] ) );
  DFFASX1 \R_reg[7][21]  ( .D(n4003), .CLK(clk), .SETB(reset_n), .Q(\R[7][21] ) );
  DFFASX1 \R_reg[7][20]  ( .D(n4002), .CLK(clk), .SETB(reset_n), .Q(\R[7][20] ) );
  DFFASX1 \R_reg[7][19]  ( .D(n4001), .CLK(clk), .SETB(reset_n), .Q(\R[7][19] ) );
  DFFASX1 \R_reg[7][18]  ( .D(n4000), .CLK(clk), .SETB(reset_n), .Q(\R[7][18] ) );
  DFFASX1 \R_reg[7][17]  ( .D(n3999), .CLK(clk), .SETB(reset_n), .Q(\R[7][17] ) );
  DFFASX1 \R_reg[7][16]  ( .D(n3998), .CLK(clk), .SETB(reset_n), .Q(\R[7][16] ) );
  DFFASX1 \R_reg[7][15]  ( .D(n3997), .CLK(clk), .SETB(reset_n), .Q(\R[7][15] ) );
  DFFASX1 \R_reg[7][14]  ( .D(n3996), .CLK(clk), .SETB(reset_n), .Q(\R[7][14] ) );
  DFFASX1 \R_reg[7][13]  ( .D(n3995), .CLK(clk), .SETB(reset_n), .Q(\R[7][13] ) );
  DFFASX1 \R_reg[7][12]  ( .D(n3994), .CLK(clk), .SETB(reset_n), .Q(\R[7][12] ) );
  DFFASX1 \R_reg[7][11]  ( .D(n3993), .CLK(clk), .SETB(reset_n), .Q(\R[7][11] ) );
  DFFASX1 \R_reg[7][10]  ( .D(n3992), .CLK(clk), .SETB(reset_n), .Q(\R[7][10] ) );
  DFFASX1 \R_reg[7][9]  ( .D(n3991), .CLK(clk), .SETB(reset_n), .Q(\R[7][9] )
         );
  DFFASX1 \R_reg[7][8]  ( .D(n3990), .CLK(clk), .SETB(reset_n), .Q(\R[7][8] )
         );
  DFFASX1 \R_reg[7][7]  ( .D(n3989), .CLK(clk), .SETB(reset_n), .Q(\R[7][7] )
         );
  DFFASX1 \R_reg[7][6]  ( .D(n3988), .CLK(clk), .SETB(reset_n), .Q(\R[7][6] )
         );
  DFFASX1 \R_reg[7][5]  ( .D(n3987), .CLK(clk), .SETB(reset_n), .Q(\R[7][5] )
         );
  DFFASX1 \R_reg[7][4]  ( .D(n3986), .CLK(clk), .SETB(reset_n), .Q(\R[7][4] )
         );
  DFFASX1 \R_reg[7][3]  ( .D(n3985), .CLK(clk), .SETB(reset_n), .Q(\R[7][3] )
         );
  DFFASX1 \R_reg[7][2]  ( .D(n3984), .CLK(clk), .SETB(reset_n), .Q(\R[7][2] )
         );
  DFFASX1 \R_reg[7][1]  ( .D(n3983), .CLK(clk), .SETB(reset_n), .Q(\R[7][1] )
         );
  DFFASX1 \R_reg[7][0]  ( .D(n3982), .CLK(clk), .SETB(reset_n), .Q(\R[7][0] )
         );
  DFFASX1 \R_reg[6][31]  ( .D(n3981), .CLK(clk), .SETB(reset_n), .Q(\R[6][31] ) );
  DFFASX1 \R_reg[6][30]  ( .D(n3980), .CLK(clk), .SETB(reset_n), .Q(\R[6][30] ) );
  DFFASX1 \R_reg[6][29]  ( .D(n3979), .CLK(clk), .SETB(reset_n), .Q(\R[6][29] ) );
  DFFASX1 \R_reg[6][28]  ( .D(n3978), .CLK(clk), .SETB(reset_n), .Q(\R[6][28] ) );
  DFFASX1 \R_reg[6][27]  ( .D(n3977), .CLK(clk), .SETB(reset_n), .Q(\R[6][27] ) );
  DFFASX1 \R_reg[6][26]  ( .D(n3976), .CLK(clk), .SETB(reset_n), .Q(\R[6][26] ) );
  DFFASX1 \R_reg[6][25]  ( .D(n3975), .CLK(clk), .SETB(reset_n), .Q(\R[6][25] ) );
  DFFASX1 \R_reg[6][24]  ( .D(n3974), .CLK(clk), .SETB(reset_n), .Q(\R[6][24] ) );
  DFFASX1 \R_reg[6][23]  ( .D(n3973), .CLK(clk), .SETB(reset_n), .Q(\R[6][23] ) );
  DFFASX1 \R_reg[6][22]  ( .D(n3972), .CLK(clk), .SETB(reset_n), .Q(\R[6][22] ) );
  DFFASX1 \R_reg[6][21]  ( .D(n3971), .CLK(clk), .SETB(reset_n), .Q(\R[6][21] ) );
  DFFASX1 \R_reg[6][20]  ( .D(n3970), .CLK(clk), .SETB(reset_n), .Q(\R[6][20] ) );
  DFFASX1 \R_reg[6][19]  ( .D(n3969), .CLK(clk), .SETB(reset_n), .Q(\R[6][19] ) );
  DFFASX1 \R_reg[6][18]  ( .D(n3968), .CLK(clk), .SETB(reset_n), .Q(\R[6][18] ) );
  DFFASX1 \R_reg[6][17]  ( .D(n3967), .CLK(clk), .SETB(reset_n), .Q(\R[6][17] ) );
  DFFASX1 \R_reg[6][16]  ( .D(n3966), .CLK(clk), .SETB(reset_n), .Q(\R[6][16] ) );
  DFFASX1 \R_reg[6][15]  ( .D(n3965), .CLK(clk), .SETB(reset_n), .Q(\R[6][15] ) );
  DFFASX1 \R_reg[6][14]  ( .D(n3964), .CLK(clk), .SETB(reset_n), .Q(\R[6][14] ) );
  DFFASX1 \R_reg[6][13]  ( .D(n3963), .CLK(clk), .SETB(reset_n), .Q(\R[6][13] ) );
  DFFASX1 \R_reg[6][12]  ( .D(n3962), .CLK(clk), .SETB(reset_n), .Q(\R[6][12] ) );
  DFFASX1 \R_reg[6][11]  ( .D(n3961), .CLK(clk), .SETB(reset_n), .Q(\R[6][11] ) );
  DFFASX1 \R_reg[6][10]  ( .D(n3960), .CLK(clk), .SETB(reset_n), .Q(\R[6][10] ) );
  DFFASX1 \R_reg[6][9]  ( .D(n3959), .CLK(clk), .SETB(reset_n), .Q(\R[6][9] )
         );
  DFFASX1 \R_reg[6][8]  ( .D(n3958), .CLK(clk), .SETB(reset_n), .Q(\R[6][8] )
         );
  DFFASX1 \R_reg[6][7]  ( .D(n3957), .CLK(clk), .SETB(reset_n), .Q(\R[6][7] )
         );
  DFFASX1 \R_reg[6][6]  ( .D(n3956), .CLK(clk), .SETB(reset_n), .Q(\R[6][6] )
         );
  DFFASX1 \R_reg[6][5]  ( .D(n3955), .CLK(clk), .SETB(reset_n), .Q(\R[6][5] )
         );
  DFFASX1 \R_reg[6][4]  ( .D(n3954), .CLK(clk), .SETB(reset_n), .Q(\R[6][4] )
         );
  DFFASX1 \R_reg[6][3]  ( .D(n3953), .CLK(clk), .SETB(reset_n), .Q(\R[6][3] )
         );
  DFFASX1 \R_reg[6][2]  ( .D(n3952), .CLK(clk), .SETB(reset_n), .Q(\R[6][2] )
         );
  DFFASX1 \R_reg[6][1]  ( .D(n3951), .CLK(clk), .SETB(reset_n), .Q(\R[6][1] )
         );
  DFFASX1 \R_reg[6][0]  ( .D(n3950), .CLK(clk), .SETB(reset_n), .Q(\R[6][0] )
         );
  DFFASX1 \R_reg[5][31]  ( .D(n3949), .CLK(clk), .SETB(reset_n), .Q(\R[5][31] ) );
  DFFASX1 \R_reg[5][30]  ( .D(n3948), .CLK(clk), .SETB(reset_n), .Q(\R[5][30] ) );
  DFFASX1 \R_reg[5][29]  ( .D(n3947), .CLK(clk), .SETB(reset_n), .Q(\R[5][29] ) );
  DFFASX1 \R_reg[5][28]  ( .D(n3946), .CLK(clk), .SETB(reset_n), .Q(\R[5][28] ) );
  DFFASX1 \R_reg[5][27]  ( .D(n3945), .CLK(clk), .SETB(reset_n), .Q(\R[5][27] ) );
  DFFASX1 \R_reg[5][26]  ( .D(n3944), .CLK(clk), .SETB(reset_n), .Q(\R[5][26] ) );
  DFFASX1 \R_reg[5][25]  ( .D(n3943), .CLK(clk), .SETB(reset_n), .Q(\R[5][25] ) );
  DFFASX1 \R_reg[5][24]  ( .D(n3942), .CLK(clk), .SETB(reset_n), .Q(\R[5][24] ) );
  DFFASX1 \R_reg[5][23]  ( .D(n3941), .CLK(clk), .SETB(reset_n), .Q(\R[5][23] ) );
  DFFASX1 \R_reg[5][22]  ( .D(n3940), .CLK(clk), .SETB(reset_n), .Q(\R[5][22] ) );
  DFFASX1 \R_reg[5][21]  ( .D(n3939), .CLK(clk), .SETB(reset_n), .Q(\R[5][21] ) );
  DFFASX1 \R_reg[5][20]  ( .D(n3938), .CLK(clk), .SETB(reset_n), .Q(\R[5][20] ) );
  DFFASX1 \R_reg[5][19]  ( .D(n3937), .CLK(clk), .SETB(reset_n), .Q(\R[5][19] ) );
  DFFASX1 \R_reg[5][18]  ( .D(n3936), .CLK(clk), .SETB(reset_n), .Q(\R[5][18] ) );
  DFFASX1 \R_reg[5][17]  ( .D(n3935), .CLK(clk), .SETB(reset_n), .Q(\R[5][17] ) );
  DFFASX1 \R_reg[5][16]  ( .D(n3934), .CLK(clk), .SETB(reset_n), .Q(\R[5][16] ) );
  DFFASX1 \R_reg[5][15]  ( .D(n3933), .CLK(clk), .SETB(reset_n), .Q(\R[5][15] ) );
  DFFASX1 \R_reg[5][14]  ( .D(n3932), .CLK(clk), .SETB(reset_n), .Q(\R[5][14] ) );
  DFFASX1 \R_reg[5][13]  ( .D(n3931), .CLK(clk), .SETB(reset_n), .Q(\R[5][13] ) );
  DFFASX1 \R_reg[5][12]  ( .D(n3930), .CLK(clk), .SETB(reset_n), .Q(\R[5][12] ) );
  DFFASX1 \R_reg[5][11]  ( .D(n3929), .CLK(clk), .SETB(reset_n), .Q(\R[5][11] ) );
  DFFASX1 \R_reg[5][10]  ( .D(n3928), .CLK(clk), .SETB(reset_n), .Q(\R[5][10] ) );
  DFFASX1 \R_reg[5][9]  ( .D(n3927), .CLK(clk), .SETB(reset_n), .Q(\R[5][9] )
         );
  DFFASX1 \R_reg[5][8]  ( .D(n3926), .CLK(clk), .SETB(reset_n), .Q(\R[5][8] )
         );
  DFFASX1 \R_reg[5][7]  ( .D(n3925), .CLK(clk), .SETB(reset_n), .Q(\R[5][7] )
         );
  DFFASX1 \R_reg[5][6]  ( .D(n3924), .CLK(clk), .SETB(reset_n), .Q(\R[5][6] )
         );
  DFFASX1 \R_reg[5][5]  ( .D(n3923), .CLK(clk), .SETB(reset_n), .Q(\R[5][5] )
         );
  DFFASX1 \R_reg[5][4]  ( .D(n3922), .CLK(clk), .SETB(reset_n), .Q(\R[5][4] )
         );
  DFFASX1 \R_reg[5][3]  ( .D(n3921), .CLK(clk), .SETB(reset_n), .Q(\R[5][3] )
         );
  DFFASX1 \R_reg[5][2]  ( .D(n3920), .CLK(clk), .SETB(reset_n), .Q(\R[5][2] )
         );
  DFFASX1 \R_reg[5][1]  ( .D(n3919), .CLK(clk), .SETB(reset_n), .Q(\R[5][1] )
         );
  DFFASX1 \R_reg[5][0]  ( .D(n3918), .CLK(clk), .SETB(reset_n), .Q(\R[5][0] )
         );
  DFFASX1 \R_reg[4][31]  ( .D(n3917), .CLK(clk), .SETB(reset_n), .Q(\R[4][31] ) );
  DFFASX1 \R_reg[4][30]  ( .D(n3916), .CLK(clk), .SETB(reset_n), .Q(\R[4][30] ) );
  DFFASX1 \R_reg[4][29]  ( .D(n3915), .CLK(clk), .SETB(reset_n), .Q(\R[4][29] ) );
  DFFASX1 \R_reg[4][28]  ( .D(n3914), .CLK(clk), .SETB(reset_n), .Q(\R[4][28] ) );
  DFFASX1 \R_reg[4][27]  ( .D(n3913), .CLK(clk), .SETB(reset_n), .Q(\R[4][27] ) );
  DFFASX1 \R_reg[4][26]  ( .D(n3912), .CLK(clk), .SETB(reset_n), .Q(\R[4][26] ) );
  DFFASX1 \R_reg[4][25]  ( .D(n3911), .CLK(clk), .SETB(reset_n), .Q(\R[4][25] ) );
  DFFASX1 \R_reg[4][24]  ( .D(n3910), .CLK(clk), .SETB(reset_n), .Q(\R[4][24] ) );
  DFFASX1 \R_reg[4][23]  ( .D(n3909), .CLK(clk), .SETB(reset_n), .Q(\R[4][23] ) );
  DFFASX1 \R_reg[4][22]  ( .D(n3908), .CLK(clk), .SETB(reset_n), .Q(\R[4][22] ) );
  DFFASX1 \R_reg[4][21]  ( .D(n3907), .CLK(clk), .SETB(reset_n), .Q(\R[4][21] ) );
  DFFASX1 \R_reg[4][20]  ( .D(n3906), .CLK(clk), .SETB(reset_n), .Q(\R[4][20] ) );
  DFFASX1 \R_reg[4][19]  ( .D(n3905), .CLK(clk), .SETB(reset_n), .Q(\R[4][19] ) );
  DFFASX1 \R_reg[4][18]  ( .D(n3904), .CLK(clk), .SETB(reset_n), .Q(\R[4][18] ) );
  DFFASX1 \R_reg[4][17]  ( .D(n3903), .CLK(clk), .SETB(reset_n), .Q(\R[4][17] ) );
  DFFASX1 \R_reg[4][16]  ( .D(n3902), .CLK(clk), .SETB(reset_n), .Q(\R[4][16] ) );
  DFFASX1 \R_reg[4][15]  ( .D(n3901), .CLK(clk), .SETB(reset_n), .Q(\R[4][15] ) );
  DFFASX1 \R_reg[4][14]  ( .D(n3900), .CLK(clk), .SETB(reset_n), .Q(\R[4][14] ) );
  DFFASX1 \R_reg[4][13]  ( .D(n3899), .CLK(clk), .SETB(reset_n), .Q(\R[4][13] ) );
  DFFASX1 \R_reg[4][12]  ( .D(n3898), .CLK(clk), .SETB(reset_n), .Q(\R[4][12] ) );
  DFFASX1 \R_reg[4][11]  ( .D(n3897), .CLK(clk), .SETB(reset_n), .Q(\R[4][11] ) );
  DFFASX1 \R_reg[4][10]  ( .D(n3896), .CLK(clk), .SETB(reset_n), .Q(\R[4][10] ) );
  DFFASX1 \R_reg[4][9]  ( .D(n3895), .CLK(clk), .SETB(reset_n), .Q(\R[4][9] )
         );
  DFFASX1 \R_reg[4][8]  ( .D(n3894), .CLK(clk), .SETB(reset_n), .Q(\R[4][8] )
         );
  DFFASX1 \R_reg[4][7]  ( .D(n3893), .CLK(clk), .SETB(reset_n), .Q(\R[4][7] )
         );
  DFFASX1 \R_reg[4][6]  ( .D(n3892), .CLK(clk), .SETB(reset_n), .Q(\R[4][6] )
         );
  DFFASX1 \R_reg[4][5]  ( .D(n3891), .CLK(clk), .SETB(reset_n), .Q(\R[4][5] )
         );
  DFFASX1 \R_reg[4][4]  ( .D(n3890), .CLK(clk), .SETB(reset_n), .Q(\R[4][4] )
         );
  DFFASX1 \R_reg[4][3]  ( .D(n3889), .CLK(clk), .SETB(reset_n), .Q(\R[4][3] )
         );
  DFFASX1 \R_reg[4][2]  ( .D(n3888), .CLK(clk), .SETB(reset_n), .Q(\R[4][2] )
         );
  DFFASX1 \R_reg[4][1]  ( .D(n3887), .CLK(clk), .SETB(reset_n), .Q(\R[4][1] )
         );
  DFFASX1 \R_reg[4][0]  ( .D(n3886), .CLK(clk), .SETB(reset_n), .Q(\R[4][0] )
         );
  DFFASX1 \R_reg[3][31]  ( .D(n3885), .CLK(clk), .SETB(reset_n), .Q(\R[3][31] ) );
  DFFASX1 \R_reg[3][30]  ( .D(n3884), .CLK(clk), .SETB(reset_n), .Q(\R[3][30] ) );
  DFFASX1 \R_reg[3][29]  ( .D(n3883), .CLK(clk), .SETB(reset_n), .Q(\R[3][29] ) );
  DFFASX1 \R_reg[3][28]  ( .D(n3882), .CLK(clk), .SETB(reset_n), .Q(\R[3][28] ) );
  DFFASX1 \R_reg[3][27]  ( .D(n3881), .CLK(clk), .SETB(reset_n), .Q(\R[3][27] ) );
  DFFASX1 \R_reg[3][26]  ( .D(n3880), .CLK(clk), .SETB(reset_n), .Q(\R[3][26] ) );
  DFFASX1 \R_reg[3][25]  ( .D(n3879), .CLK(clk), .SETB(reset_n), .Q(\R[3][25] ) );
  DFFASX1 \R_reg[3][24]  ( .D(n3878), .CLK(clk), .SETB(reset_n), .Q(\R[3][24] ) );
  DFFASX1 \R_reg[3][23]  ( .D(n3877), .CLK(clk), .SETB(reset_n), .Q(\R[3][23] ) );
  DFFASX1 \R_reg[3][22]  ( .D(n3876), .CLK(clk), .SETB(reset_n), .Q(\R[3][22] ) );
  DFFASX1 \R_reg[3][21]  ( .D(n3875), .CLK(clk), .SETB(reset_n), .Q(\R[3][21] ) );
  DFFASX1 \R_reg[3][20]  ( .D(n3874), .CLK(clk), .SETB(reset_n), .Q(\R[3][20] ) );
  DFFASX1 \R_reg[3][19]  ( .D(n3873), .CLK(clk), .SETB(reset_n), .Q(\R[3][19] ) );
  DFFASX1 \R_reg[3][18]  ( .D(n3872), .CLK(clk), .SETB(reset_n), .Q(\R[3][18] ) );
  DFFASX1 \R_reg[3][17]  ( .D(n3871), .CLK(clk), .SETB(reset_n), .Q(\R[3][17] ) );
  DFFASX1 \R_reg[3][16]  ( .D(n3870), .CLK(clk), .SETB(reset_n), .Q(\R[3][16] ) );
  DFFASX1 \R_reg[3][15]  ( .D(n3869), .CLK(clk), .SETB(reset_n), .Q(\R[3][15] ) );
  DFFASX1 \R_reg[3][14]  ( .D(n3868), .CLK(clk), .SETB(reset_n), .Q(\R[3][14] ) );
  DFFASX1 \R_reg[3][13]  ( .D(n3867), .CLK(clk), .SETB(reset_n), .Q(\R[3][13] ) );
  DFFASX1 \R_reg[3][12]  ( .D(n3866), .CLK(clk), .SETB(reset_n), .Q(\R[3][12] ) );
  DFFASX1 \R_reg[3][11]  ( .D(n3865), .CLK(clk), .SETB(reset_n), .Q(\R[3][11] ) );
  DFFASX1 \R_reg[3][10]  ( .D(n3864), .CLK(clk), .SETB(reset_n), .Q(\R[3][10] ) );
  DFFASX1 \R_reg[3][9]  ( .D(n3863), .CLK(clk), .SETB(reset_n), .Q(\R[3][9] )
         );
  DFFASX1 \R_reg[3][8]  ( .D(n3862), .CLK(clk), .SETB(reset_n), .Q(\R[3][8] )
         );
  DFFASX1 \R_reg[3][7]  ( .D(n3861), .CLK(clk), .SETB(reset_n), .Q(\R[3][7] )
         );
  DFFASX1 \R_reg[3][6]  ( .D(n3860), .CLK(clk), .SETB(reset_n), .Q(\R[3][6] )
         );
  DFFASX1 \R_reg[3][5]  ( .D(n3859), .CLK(clk), .SETB(reset_n), .Q(\R[3][5] )
         );
  DFFASX1 \R_reg[3][4]  ( .D(n3858), .CLK(clk), .SETB(reset_n), .Q(\R[3][4] )
         );
  DFFASX1 \R_reg[3][3]  ( .D(n3857), .CLK(clk), .SETB(reset_n), .Q(\R[3][3] )
         );
  DFFASX1 \R_reg[3][2]  ( .D(n3856), .CLK(clk), .SETB(reset_n), .Q(\R[3][2] )
         );
  DFFASX1 \R_reg[3][1]  ( .D(n3855), .CLK(clk), .SETB(reset_n), .Q(\R[3][1] )
         );
  DFFASX1 \R_reg[3][0]  ( .D(n3854), .CLK(clk), .SETB(reset_n), .Q(\R[3][0] )
         );
  DFFASX1 \R_reg[2][31]  ( .D(n3853), .CLK(clk), .SETB(reset_n), .Q(\R[2][31] ) );
  DFFASX1 \R_reg[2][30]  ( .D(n3852), .CLK(clk), .SETB(reset_n), .Q(\R[2][30] ) );
  DFFASX1 \R_reg[2][29]  ( .D(n3851), .CLK(clk), .SETB(reset_n), .Q(\R[2][29] ) );
  DFFASX1 \R_reg[2][28]  ( .D(n3850), .CLK(clk), .SETB(reset_n), .Q(\R[2][28] ) );
  DFFASX1 \R_reg[2][27]  ( .D(n3849), .CLK(clk), .SETB(reset_n), .Q(\R[2][27] ) );
  DFFASX1 \R_reg[2][26]  ( .D(n3848), .CLK(clk), .SETB(reset_n), .Q(\R[2][26] ) );
  DFFASX1 \R_reg[2][25]  ( .D(n3847), .CLK(clk), .SETB(reset_n), .Q(\R[2][25] ) );
  DFFASX1 \R_reg[2][24]  ( .D(n3846), .CLK(clk), .SETB(reset_n), .Q(\R[2][24] ) );
  DFFASX1 \R_reg[2][23]  ( .D(n3845), .CLK(clk), .SETB(reset_n), .Q(\R[2][23] ) );
  DFFASX1 \R_reg[2][22]  ( .D(n3844), .CLK(clk), .SETB(reset_n), .Q(\R[2][22] ) );
  DFFASX1 \R_reg[2][21]  ( .D(n3843), .CLK(clk), .SETB(reset_n), .Q(\R[2][21] ) );
  DFFASX1 \R_reg[2][20]  ( .D(n3842), .CLK(clk), .SETB(reset_n), .Q(\R[2][20] ) );
  DFFASX1 \R_reg[2][19]  ( .D(n3841), .CLK(clk), .SETB(reset_n), .Q(\R[2][19] ) );
  DFFASX1 \R_reg[2][18]  ( .D(n3840), .CLK(clk), .SETB(reset_n), .Q(\R[2][18] ) );
  DFFASX1 \R_reg[2][17]  ( .D(n3839), .CLK(clk), .SETB(reset_n), .Q(\R[2][17] ) );
  DFFASX1 \R_reg[2][16]  ( .D(n3838), .CLK(clk), .SETB(reset_n), .Q(\R[2][16] ) );
  DFFASX1 \R_reg[2][15]  ( .D(n3837), .CLK(clk), .SETB(reset_n), .Q(\R[2][15] ) );
  DFFASX1 \R_reg[2][14]  ( .D(n3836), .CLK(clk), .SETB(reset_n), .Q(\R[2][14] ) );
  DFFASX1 \R_reg[2][13]  ( .D(n3835), .CLK(clk), .SETB(reset_n), .Q(\R[2][13] ) );
  DFFASX1 \R_reg[2][12]  ( .D(n3834), .CLK(clk), .SETB(reset_n), .Q(\R[2][12] ) );
  DFFASX1 \R_reg[2][11]  ( .D(n3833), .CLK(clk), .SETB(reset_n), .Q(\R[2][11] ) );
  DFFASX1 \R_reg[2][10]  ( .D(n3832), .CLK(clk), .SETB(reset_n), .Q(\R[2][10] ) );
  DFFASX1 \R_reg[2][9]  ( .D(n3831), .CLK(clk), .SETB(reset_n), .Q(\R[2][9] )
         );
  DFFASX1 \R_reg[2][8]  ( .D(n3830), .CLK(clk), .SETB(reset_n), .Q(\R[2][8] )
         );
  DFFASX1 \R_reg[2][7]  ( .D(n3829), .CLK(clk), .SETB(reset_n), .Q(\R[2][7] )
         );
  DFFASX1 \R_reg[2][6]  ( .D(n3828), .CLK(clk), .SETB(reset_n), .Q(\R[2][6] )
         );
  DFFASX1 \R_reg[2][5]  ( .D(n3827), .CLK(clk), .SETB(reset_n), .Q(\R[2][5] )
         );
  DFFASX1 \R_reg[2][4]  ( .D(n3826), .CLK(clk), .SETB(reset_n), .Q(\R[2][4] )
         );
  DFFASX1 \R_reg[2][3]  ( .D(n3825), .CLK(clk), .SETB(reset_n), .Q(\R[2][3] )
         );
  DFFASX1 \R_reg[2][2]  ( .D(n3824), .CLK(clk), .SETB(reset_n), .Q(\R[2][2] )
         );
  DFFASX1 \R_reg[2][1]  ( .D(n3823), .CLK(clk), .SETB(reset_n), .Q(\R[2][1] )
         );
  DFFASX1 \R_reg[2][0]  ( .D(n3822), .CLK(clk), .SETB(reset_n), .Q(\R[2][0] )
         );
  DFFASX1 \R_reg[1][31]  ( .D(n3821), .CLK(clk), .SETB(reset_n), .Q(\R[1][31] ) );
  DFFASX1 \R_reg[1][30]  ( .D(n3820), .CLK(clk), .SETB(reset_n), .Q(\R[1][30] ) );
  DFFASX1 \R_reg[1][29]  ( .D(n3819), .CLK(clk), .SETB(reset_n), .Q(\R[1][29] ) );
  DFFASX1 \R_reg[1][28]  ( .D(n3818), .CLK(clk), .SETB(reset_n), .Q(\R[1][28] ) );
  DFFASX1 \R_reg[1][27]  ( .D(n3817), .CLK(clk), .SETB(reset_n), .Q(\R[1][27] ) );
  DFFASX1 \R_reg[1][26]  ( .D(n3816), .CLK(clk), .SETB(reset_n), .Q(\R[1][26] ) );
  DFFASX1 \R_reg[1][25]  ( .D(n3815), .CLK(clk), .SETB(reset_n), .Q(\R[1][25] ) );
  DFFASX1 \R_reg[1][24]  ( .D(n3814), .CLK(clk), .SETB(reset_n), .Q(\R[1][24] ) );
  DFFASX1 \R_reg[1][23]  ( .D(n3813), .CLK(clk), .SETB(reset_n), .Q(\R[1][23] ) );
  DFFASX1 \R_reg[1][22]  ( .D(n3812), .CLK(clk), .SETB(reset_n), .Q(\R[1][22] ) );
  DFFASX1 \R_reg[1][21]  ( .D(n3811), .CLK(clk), .SETB(reset_n), .Q(\R[1][21] ) );
  DFFASX1 \R_reg[1][20]  ( .D(n3810), .CLK(clk), .SETB(reset_n), .Q(\R[1][20] ) );
  DFFASX1 \R_reg[1][19]  ( .D(n3809), .CLK(clk), .SETB(reset_n), .Q(\R[1][19] ) );
  DFFASX1 \R_reg[1][18]  ( .D(n3808), .CLK(clk), .SETB(reset_n), .Q(\R[1][18] ) );
  DFFASX1 \R_reg[1][17]  ( .D(n3807), .CLK(clk), .SETB(reset_n), .Q(\R[1][17] ) );
  DFFASX1 \R_reg[1][16]  ( .D(n3806), .CLK(clk), .SETB(reset_n), .Q(\R[1][16] ) );
  DFFASX1 \R_reg[1][15]  ( .D(n3805), .CLK(clk), .SETB(reset_n), .Q(\R[1][15] ) );
  DFFASX1 \R_reg[1][14]  ( .D(n3804), .CLK(clk), .SETB(reset_n), .Q(\R[1][14] ) );
  DFFASX1 \R_reg[1][13]  ( .D(n3803), .CLK(clk), .SETB(reset_n), .Q(\R[1][13] ) );
  DFFASX1 \R_reg[1][12]  ( .D(n3802), .CLK(clk), .SETB(reset_n), .Q(\R[1][12] ) );
  DFFASX1 \R_reg[1][11]  ( .D(n3801), .CLK(clk), .SETB(reset_n), .Q(\R[1][11] ) );
  DFFASX1 \R_reg[1][10]  ( .D(n3800), .CLK(clk), .SETB(reset_n), .Q(\R[1][10] ) );
  DFFASX1 \R_reg[1][9]  ( .D(n3799), .CLK(clk), .SETB(reset_n), .Q(\R[1][9] )
         );
  DFFASX1 \R_reg[1][8]  ( .D(n3798), .CLK(clk), .SETB(reset_n), .Q(\R[1][8] )
         );
  DFFASX1 \R_reg[1][7]  ( .D(n3797), .CLK(clk), .SETB(reset_n), .Q(\R[1][7] )
         );
  DFFASX1 \R_reg[1][6]  ( .D(n3796), .CLK(clk), .SETB(reset_n), .Q(\R[1][6] )
         );
  DFFASX1 \R_reg[1][5]  ( .D(n3795), .CLK(clk), .SETB(reset_n), .Q(\R[1][5] )
         );
  DFFASX1 \R_reg[1][4]  ( .D(n3794), .CLK(clk), .SETB(reset_n), .Q(\R[1][4] )
         );
  DFFASX1 \R_reg[1][3]  ( .D(n3793), .CLK(clk), .SETB(reset_n), .Q(\R[1][3] )
         );
  DFFASX1 \R_reg[1][2]  ( .D(n3792), .CLK(clk), .SETB(reset_n), .Q(\R[1][2] )
         );
  DFFASX1 \R_reg[1][1]  ( .D(n3791), .CLK(clk), .SETB(reset_n), .Q(\R[1][1] )
         );
  DFFASX1 \R_reg[1][0]  ( .D(n3790), .CLK(clk), .SETB(reset_n), .Q(\R[1][0] )
         );
  DFFASX1 \R_reg[0][31]  ( .D(n3789), .CLK(clk), .SETB(reset_n), .Q(\R[0][31] ) );
  DFFASX1 \R_reg[0][30]  ( .D(n3788), .CLK(clk), .SETB(reset_n), .Q(\R[0][30] ) );
  DFFASX1 \R_reg[0][29]  ( .D(n3787), .CLK(clk), .SETB(reset_n), .Q(\R[0][29] ) );
  DFFASX1 \R_reg[0][28]  ( .D(n3786), .CLK(clk), .SETB(reset_n), .Q(\R[0][28] ) );
  DFFASX1 \R_reg[0][27]  ( .D(n3785), .CLK(clk), .SETB(reset_n), .Q(\R[0][27] ) );
  DFFASX1 \R_reg[0][26]  ( .D(n3784), .CLK(clk), .SETB(reset_n), .Q(\R[0][26] ) );
  DFFASX1 \R_reg[0][25]  ( .D(n3783), .CLK(clk), .SETB(reset_n), .Q(\R[0][25] ) );
  DFFASX1 \R_reg[0][24]  ( .D(n3782), .CLK(clk), .SETB(reset_n), .Q(\R[0][24] ) );
  DFFASX1 \R_reg[0][23]  ( .D(n3781), .CLK(clk), .SETB(reset_n), .Q(\R[0][23] ) );
  DFFASX1 \R_reg[0][22]  ( .D(n3780), .CLK(clk), .SETB(reset_n), .Q(\R[0][22] ) );
  DFFASX1 \R_reg[0][21]  ( .D(n3779), .CLK(clk), .SETB(reset_n), .Q(\R[0][21] ) );
  DFFASX1 \R_reg[0][20]  ( .D(n3778), .CLK(clk), .SETB(reset_n), .Q(\R[0][20] ) );
  DFFASX1 \R_reg[0][19]  ( .D(n3777), .CLK(clk), .SETB(reset_n), .Q(\R[0][19] ) );
  DFFASX1 \R_reg[0][18]  ( .D(n3776), .CLK(clk), .SETB(reset_n), .Q(\R[0][18] ) );
  DFFASX1 \R_reg[0][17]  ( .D(n3775), .CLK(clk), .SETB(reset_n), .Q(\R[0][17] ) );
  DFFASX1 \R_reg[0][16]  ( .D(n3774), .CLK(clk), .SETB(reset_n), .Q(\R[0][16] ) );
  DFFASX1 \R_reg[0][15]  ( .D(n3773), .CLK(clk), .SETB(reset_n), .Q(\R[0][15] ) );
  DFFASX1 \R_reg[0][14]  ( .D(n3772), .CLK(clk), .SETB(reset_n), .Q(\R[0][14] ) );
  DFFASX1 \R_reg[0][13]  ( .D(n3771), .CLK(clk), .SETB(reset_n), .Q(\R[0][13] ) );
  DFFASX1 \R_reg[0][12]  ( .D(n3770), .CLK(clk), .SETB(reset_n), .Q(\R[0][12] ) );
  DFFASX1 \R_reg[0][11]  ( .D(n3769), .CLK(clk), .SETB(reset_n), .Q(\R[0][11] ) );
  DFFASX1 \R_reg[0][10]  ( .D(n3768), .CLK(clk), .SETB(reset_n), .Q(\R[0][10] ) );
  DFFASX1 \R_reg[0][9]  ( .D(n3767), .CLK(clk), .SETB(reset_n), .Q(\R[0][9] )
         );
  DFFASX1 \R_reg[0][8]  ( .D(n3766), .CLK(clk), .SETB(reset_n), .Q(\R[0][8] )
         );
  DFFASX1 \R_reg[0][7]  ( .D(n3765), .CLK(clk), .SETB(reset_n), .Q(\R[0][7] )
         );
  DFFASX1 \R_reg[0][6]  ( .D(n3764), .CLK(clk), .SETB(reset_n), .Q(\R[0][6] )
         );
  DFFASX1 \R_reg[0][5]  ( .D(n3763), .CLK(clk), .SETB(reset_n), .Q(\R[0][5] )
         );
  DFFASX1 \R_reg[0][4]  ( .D(n3762), .CLK(clk), .SETB(reset_n), .Q(\R[0][4] )
         );
  DFFASX1 \R_reg[0][3]  ( .D(n3761), .CLK(clk), .SETB(reset_n), .Q(\R[0][3] )
         );
  DFFASX1 \R_reg[0][2]  ( .D(n3760), .CLK(clk), .SETB(reset_n), .Q(\R[0][2] )
         );
  DFFASX1 \R_reg[0][1]  ( .D(n3759), .CLK(clk), .SETB(reset_n), .Q(\R[0][1] )
         );
  DFFASX1 \R_reg[0][0]  ( .D(n3758), .CLK(clk), .SETB(reset_n), .Q(\R[0][0] )
         );
  thumb_DW01_addsub_0 sub_0_root_sub_760_2 ( .A({n393, n394, n395, n396, n397, 
        n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
        n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
        n422, n423, n424, n425}), .B({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, n4486}), .CI(1'b0), .ADD_SUB(1'b1), .SUM({N5292, N5291, N5290, 
        N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, 
        N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, 
        N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260})
         );
  thumb_DW01_addsub_1 r1728 ( .A({1'b0, \U3/U87/Z_31 , \U3/U87/Z_30 , 
        \U3/U87/Z_29 , \U3/U87/Z_28 , \U3/U87/Z_27 , \U3/U87/Z_26 , 
        \U3/U87/Z_25 , \U3/U87/Z_24 , \U3/U87/Z_23 , \U3/U87/Z_22 , 
        \U3/U87/Z_21 , \U3/U87/Z_20 , \U3/U87/Z_19 , \U3/U87/Z_18 , 
        \U3/U87/Z_17 , \U3/U87/Z_16 , \U3/U87/Z_15 , \U3/U87/Z_14 , 
        \U3/U87/Z_13 , \U3/U87/Z_12 , \U3/U87/Z_11 , \U3/U87/Z_10 , 
        \U3/U87/Z_9 , \U3/U87/Z_8 , \U3/U87/Z_7 , \U3/U87/Z_6 , \U3/U87/Z_5 , 
        \U3/U87/Z_4 , \U3/U87/Z_3 , \U3/U87/Z_2 , \U3/U87/Z_1 , \U3/U87/Z_0 }), 
        .B({\U3/U88/Z_32 , \U3/U88/Z_31 , \U3/U88/Z_30 , \U3/U88/Z_29 , 
        \U3/U88/Z_28 , \U3/U88/Z_27 , \U3/U88/Z_26 , \U3/U88/Z_25 , 
        \U3/U88/Z_24 , \U3/U88/Z_23 , \U3/U88/Z_22 , \U3/U88/Z_21 , 
        \U3/U88/Z_20 , \U3/U88/Z_19 , \U3/U88/Z_18 , \U3/U88/Z_17 , 
        \U3/U88/Z_16 , \U3/U88/Z_15 , \U3/U88/Z_14 , \U3/U88/Z_13 , 
        \U3/U88/Z_12 , \U3/U88/Z_11 , \U3/U88/Z_10 , \U3/U88/Z_9 , 
        \U3/U88/Z_8 , \U3/U88/Z_7 , \U3/U88/Z_6 , \U3/U88/Z_5 , \U3/U88/Z_4 , 
        \U3/U88/Z_3 , \U3/U88/Z_2 , \U3/U88/Z_1 , \U3/U88/Z_0 }), .CI(
        \U3/U89/Z_0 ), .ADD_SUB(\U3/U90/Z_0 ), .SUM({n393, n394, n395, n396, 
        n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
        n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
        n421, n422, n423, n424, n425}) );
  thumb_DW01_addsub_2 r1483 ( .A({1'b0, \U3/U91/Z_31 , \U3/U91/Z_30 , 
        \U3/U91/Z_29 , \U3/U91/Z_28 , \U3/U91/Z_27 , \U3/U91/Z_26 , 
        \U3/U91/Z_25 , \U3/U91/Z_24 , \U3/U91/Z_23 , \U3/U91/Z_22 , 
        \U3/U91/Z_21 , \U3/U91/Z_20 , \U3/U91/Z_19 , \U3/U91/Z_18 , 
        \U3/U91/Z_17 , \U3/U91/Z_16 , \U3/U91/Z_15 , \U3/U91/Z_14 , 
        \U3/U91/Z_13 , \U3/U91/Z_12 , \U3/U91/Z_11 , \U3/U91/Z_10 , 
        \U3/U91/Z_9 , \U3/U91/Z_8 , \U3/U91/Z_7 , \U3/U91/Z_6 , \U3/U91/Z_5 , 
        \U3/U91/Z_4 , \U3/U91/Z_3 , \U3/U91/Z_2 , \U3/U91/Z_1 , \U3/U91/Z_0 }), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \U3/U92/Z_11 , \U3/U92/Z_10 , \U3/U92/Z_9 , \U3/U92/Z_8 , \U3/U92/Z_7 , 
        \U3/U92/Z_6 , \U3/U92/Z_5 , \U3/U92/Z_4 , \U3/U92/Z_3 , \U3/U92/Z_2 , 
        \U3/U92/Z_1 , \U3/U92/Z_0 }), .CI(1'b0), .ADD_SUB(\U3/U93/Z_0 ), .SUM(
        {n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
        n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
        n529, n530, n531, n532, n533, n534, n535, n536, n537, n538}) );
  thumb_DW01_add_0 r1223 ( .A({1'b0, ID_Rn}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        ID_imm_offset[4:0], 1'b0}), .CI(1'b0), .SUM({N4776, N4775, N4774, 
        N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, 
        N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, 
        N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744})
         );
  thumb_DW01_add_1 r1222 ( .A({1'b0, ID_Rn}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        ID_imm_offset[4:0]}), .CI(1'b0), .SUM({N4743, N4742, N4741, N4740, 
        N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, 
        N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, 
        N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711}) );
  thumb_DW01_add_2 r1221 ( .A({1'b0, ID_Rn}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        ID_imm_offset[4:0], 1'b0, 1'b0}), .CI(1'b0), .SUM({N4611, N4610, N4609, 
        N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, 
        N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, 
        N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579})
         );
  thumb_DW01_sub_0 r1220 ( .A({1'b0, ID_Rn}), .B({1'b0, N3016, ID_Rm_Rs[30:0]}), .CI(1'b0), .DIFF({N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, 
        N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, 
        N4528, N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, 
        N4518, N4517, N4516, N4515, N4514}) );
  thumb_DW01_sub_1 r1219 ( .A({1'b0, ID_Rn}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, ID_imm_offset[7:0]}), 
        .CI(1'b0), .DIFF({N4513, N4512, N4511, N4510, N4509, N4508, N4507, 
        N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, 
        N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, 
        N4486, N4485, N4484, N4483, N4482, N4481}) );
  thumb_DW01_add_3 r1148 ( .A({1'b0, SP}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, ID_imm_offset[7:0], 1'b0, 1'b0}), 
        .CI(1'b0), .SUM({N4710, N1831, N1830, N1829, N1828, N1827, N1826, 
        N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, 
        N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, 
        N1805, N1804, N1803, N1802, N1801, N1800}) );
  thumb_DW01_add_4 r1147 ( .A({1'b0, ID_PC[31:2], 1'b0, 1'b0}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        ID_imm_offset[7:0], 1'b0, 1'b0}), .CI(1'b0), .SUM({N4677, N1799, N1798, 
        N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, 
        N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, 
        N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  thumb_DW01_add_5 r1146 ( .A({1'b0, ID_Rn}), .B({1'b0, N3016, ID_Rm_Rs[30:0]}), .CI(1'b0), .SUM({N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, 
        N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, 
        N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, 
        N1739, N1738, N1737, N1736, N1735}) );
  thumb_DW01_add_6 r1142 ( .A(instruction_address), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0}), .CI(1'b0), .SUM({N354, N353, N352, N351, 
        N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, 
        N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, 
        N326, N325, N324, N323}) );
  thumb_DW_leftsh_2 sll_722 ( .A({1'b0, N4141, ID_Rd[30:0]}), .SH(
        ID_Rm_Rs[7:0]), .B({N4845, N4844, N4843, N4842, N4841, N4840, N4839, 
        N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, 
        N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, 
        N4818, N4817, N4816, N4815, N4814, N4813}) );
  thumb_DW_rightsh_3 srl_758 ( .A({N4141, ID_Rd[30:0], 1'b0}), .DATA_TC(1'b0), 
        .SH(ID_Rm_Rs[4:0]), .B({N5226, N5225, N5224, N5223, N5222, N5221, 
        N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, 
        N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, 
        N5200, N5199, N5198, N5197, N5196, N5195, N5194}) );
  thumb_DW_mult_uns_1 mult_734 ( .a({N4141, ID_Rd[30:0]}), .b({N3016, 
        ID_Rm_Rs[30:0]}), .product({SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, N5012, N5011, N5010, N5009, N5008, N5007, 
        N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, 
        N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, 
        N4986, N4985, N4984, N4983, N4982, N4981}) );
  thumb_DW_leftsh_3 sll_720 ( .A({1'b0, N3016, ID_Rm_Rs[30:0]}), .SH(
        ID_imm_offset[4:0]), .B({N4809, N4808, N4807, N4806, N4805, N4804, 
        N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, 
        N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, 
        N4783, N4782, N4781, N4780, N4779, N4778, N4777}) );
  thumb_DW_rightsh_4 srl_725 ( .A({N3016, ID_Rm_Rs[30:0], 1'b0}), .DATA_TC(
        1'b0), .SH(ID_imm_offset[4:0]), .B({N4911, N4910, N4909, N4908, N4907, 
        N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, 
        N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, 
        N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879}) );
  thumb_DW_rightsh_5 srl_728 ( .A({N4141, ID_Rd[30:0], 1'b0}), .DATA_TC(1'b0), 
        .SH(ID_Rm_Rs[7:0]), .B({N4947, N4946, N4945, N4944, N4943, N4942, 
        N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, 
        N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, 
        N4921, N4920, N4919, N4918, N4917, N4916, N4915}) );
  BSLEX1 \data_tri[0]  ( .INOUT1(n9199), .ENB(n9198), .INOUT2(data[0]) );
  BSLEX1 \data_tri[1]  ( .INOUT1(n9200), .ENB(n9198), .INOUT2(data[1]) );
  BSLEX1 \data_tri[2]  ( .INOUT1(n9201), .ENB(n9198), .INOUT2(data[2]) );
  BSLEX1 \data_tri[3]  ( .INOUT1(n9202), .ENB(n9198), .INOUT2(data[3]) );
  BSLEX1 \data_tri[4]  ( .INOUT1(n9203), .ENB(n9198), .INOUT2(data[4]) );
  BSLEX1 \data_tri[5]  ( .INOUT1(n9204), .ENB(n9198), .INOUT2(data[5]) );
  BSLEX1 \data_tri[6]  ( .INOUT1(n9205), .ENB(n9198), .INOUT2(data[6]) );
  BSLEX1 \data_tri[8]  ( .INOUT1(n9207), .ENB(n9198), .INOUT2(data[8]) );
  BSLEX1 \data_tri[9]  ( .INOUT1(n9208), .ENB(n9198), .INOUT2(data[9]) );
  BSLEX1 \data_tri[10]  ( .INOUT1(n9209), .ENB(n9198), .INOUT2(data[10]) );
  BSLEX1 \data_tri[11]  ( .INOUT1(n9210), .ENB(n9198), .INOUT2(data[11]) );
  BSLEX1 \data_tri[12]  ( .INOUT1(n9211), .ENB(n9198), .INOUT2(data[12]) );
  BSLEX1 \data_tri[13]  ( .INOUT1(n9212), .ENB(n9198), .INOUT2(data[13]) );
  BSLEX1 \data_tri[14]  ( .INOUT1(n9213), .ENB(n9198), .INOUT2(data[14]) );
  BSLEX1 \data_tri[16]  ( .INOUT1(n9215), .ENB(n9198), .INOUT2(data[16]) );
  BSLEX1 \data_tri[17]  ( .INOUT1(n9216), .ENB(n9198), .INOUT2(data[17]) );
  BSLEX1 \data_tri[18]  ( .INOUT1(n9217), .ENB(n9198), .INOUT2(data[18]) );
  BSLEX1 \data_tri[19]  ( .INOUT1(n9218), .ENB(n9198), .INOUT2(data[19]) );
  BSLEX1 \data_tri[20]  ( .INOUT1(n9219), .ENB(n9198), .INOUT2(data[20]) );
  BSLEX1 \data_tri[21]  ( .INOUT1(n9220), .ENB(n9198), .INOUT2(data[21]) );
  BSLEX1 \data_tri[22]  ( .INOUT1(n9221), .ENB(n9198), .INOUT2(data[22]) );
  BSLEX1 \data_tri[23]  ( .INOUT1(n9222), .ENB(n9198), .INOUT2(data[23]) );
  BSLEX1 \data_tri[24]  ( .INOUT1(n9223), .ENB(n9198), .INOUT2(data[24]) );
  BSLEX1 \data_tri[25]  ( .INOUT1(n9224), .ENB(n9198), .INOUT2(data[25]) );
  BSLEX1 \data_tri[26]  ( .INOUT1(n9225), .ENB(n9198), .INOUT2(data[26]) );
  BSLEX1 \data_tri[27]  ( .INOUT1(n9226), .ENB(n9198), .INOUT2(data[27]) );
  BSLEX1 \data_tri[28]  ( .INOUT1(n9227), .ENB(n9198), .INOUT2(data[28]) );
  BSLEX1 \data_tri[29]  ( .INOUT1(n9228), .ENB(n9198), .INOUT2(data[29]) );
  BSLEX1 \data_tri[30]  ( .INOUT1(n9229), .ENB(n9198), .INOUT2(data[30]) );
  BSLEX1 \data_tri[31]  ( .INOUT1(n9230), .ENB(n9198), .INOUT2(data[31]) );
  BSLEX1 \data_tri[7]  ( .INOUT1(n9206), .ENB(n9198), .INOUT2(data[7]) );
  BSLEX1 \data_tri[15]  ( .INOUT1(n9214), .ENB(n9198), .INOUT2(data[15]) );
  DFFX2 \ID_imm_offset_reg[1]  ( .D(n4293), .CLK(clk), .Q(ID_imm_offset[1]), 
        .QN(n3714) );
  DFFX2 \ID_imm_offset_reg[2]  ( .D(n4296), .CLK(clk), .Q(ID_imm_offset[2]), 
        .QN(n3715) );
  DFFX2 \ID_imm_offset_reg[0]  ( .D(n4290), .CLK(clk), .Q(ID_imm_offset[0]), 
        .QN(n3713) );
  DFFX2 \ID_Rm_Rs_reg[1]  ( .D(n4334), .CLK(clk), .Q(ID_Rm_Rs[1]), .QN(n4484)
         );
  DFFX2 \ID_Rm_Rs_reg[0]  ( .D(n4335), .CLK(clk), .Q(ID_Rm_Rs[0]), .QN(n4485)
         );
  DFFX2 \ID_imm_offset_reg[3]  ( .D(n4298), .CLK(clk), .Q(ID_imm_offset[3]), 
        .QN(n3627) );
  DFFX2 \ID_Rm_Rs_reg[2]  ( .D(n4333), .CLK(clk), .Q(ID_Rm_Rs[2]), .QN(n4483)
         );
  DFFX2 \ID_Rm_Rs_reg[3]  ( .D(n4332), .CLK(clk), .Q(ID_Rm_Rs[3]), .QN(n4482)
         );
  AND3X1 U4740 ( .IN1(n3694), .IN2(n8413), .IN3(n3696), .Q(n5706) );
  OA21X1 U4741 ( .IN1(n8415), .IN2(n7148), .IN3(n3696), .Q(n5709) );
  AND2X1 U4742 ( .IN1(n5756), .IN2(N1801), .Q(n5711) );
  AND2X1 U4743 ( .IN1(n5756), .IN2(N1800), .Q(n5712) );
  INVX0 U4744 ( .INP(n5706), .ZN(n5715) );
  INVX0 U4745 ( .INP(n5706), .ZN(n5716) );
  INVX0 U4746 ( .INP(n5706), .ZN(n5717) );
  INVX0 U4747 ( .INP(n5706), .ZN(n5718) );
  INVX0 U4748 ( .INP(n5709), .ZN(n5719) );
  INVX0 U4749 ( .INP(n5709), .ZN(n5720) );
  INVX0 U4750 ( .INP(n5709), .ZN(n5721) );
  INVX0 U4751 ( .INP(n5709), .ZN(n5722) );
  INVX2 U4752 ( .INP(n7751), .ZN(n7643) );
  NOR2X1 U4753 ( .IN1(n7097), .IN2(n7441), .QN(n7405) );
  NAND4X1 U4754 ( .IN1(n3696), .IN2(n3694), .IN3(n3629), .IN4(n3628), .QN(N318) );
  NAND3X1 U4755 ( .IN1(n8896), .IN2(n8897), .IN3(n8861), .QN(n7626) );
  NAND3X2 U4756 ( .IN1(n7800), .IN2(n7884), .IN3(n7999), .QN(\U3/U93/Z_0 ) );
  NAND2X1 U4757 ( .IN1(n7508), .IN2(n7782), .QN(\U3/U90/Z_0 ) );
  MUX21X1 U4758 ( .IN1(ID_imm_offset[7]), .IN2(ID_imm_offset[10]), .S(n5765), 
        .Q(n5723) );
  INVX0 U4759 ( .INP(n3695), .ZN(n6942) );
  INVX0 U4760 ( .INP(n3695), .ZN(n6944) );
  INVX0 U4761 ( .INP(n3695), .ZN(n6943) );
  INVX0 U4762 ( .INP(n3695), .ZN(n6946) );
  INVX0 U4763 ( .INP(n3695), .ZN(n6945) );
  INVX0 U4764 ( .INP(n3695), .ZN(n6948) );
  INVX0 U4765 ( .INP(n3695), .ZN(n6947) );
  INVX0 U4766 ( .INP(n3695), .ZN(n6950) );
  INVX0 U4767 ( .INP(n3695), .ZN(n6949) );
  NBUFFX2 U4768 ( .INP(ID_opcode[4]), .Z(n5788) );
  NBUFFX2 U4769 ( .INP(ID_opcode[4]), .Z(n5789) );
  NBUFFX2 U4770 ( .INP(ID_opcode[4]), .Z(n5791) );
  NBUFFX2 U4771 ( .INP(ID_opcode[4]), .Z(n5790) );
  NBUFFX2 U4772 ( .INP(ID_opcode[4]), .Z(n5787) );
  NBUFFX2 U4773 ( .INP(ID_opcode[4]), .Z(n5792) );
  NBUFFX2 U4774 ( .INP(ID_opcode[4]), .Z(n5794) );
  NBUFFX2 U4775 ( .INP(ID_opcode[4]), .Z(n5795) );
  NBUFFX2 U4776 ( .INP(ID_opcode[4]), .Z(n5793) );
  NBUFFX2 U4777 ( .INP(ID_opcode[4]), .Z(n5796) );
  MUX41X1 U4778 ( .IN1(\R[3][30] ), .IN3(\R[1][30] ), .IN2(\R[2][30] ), .IN4(
        \R[0][30] ), .S0(n9196), .S1(n9197), .Q(n6798) );
  MUX41X1 U4779 ( .IN1(\R[3][28] ), .IN3(\R[1][28] ), .IN2(\R[2][28] ), .IN4(
        \R[0][28] ), .S0(n9196), .S1(n9197), .Q(n6794) );
  MUX41X1 U4780 ( .IN1(\R[3][26] ), .IN3(\R[1][26] ), .IN2(\R[2][26] ), .IN4(
        \R[0][26] ), .S0(n9196), .S1(n9197), .Q(n6790) );
  MUX41X1 U4781 ( .IN1(\R[3][23] ), .IN3(\R[1][23] ), .IN2(\R[2][23] ), .IN4(
        \R[0][23] ), .S0(n9196), .S1(n9197), .Q(n6784) );
  MUX41X1 U4782 ( .IN1(\R[3][21] ), .IN3(\R[1][21] ), .IN2(\R[2][21] ), .IN4(
        \R[0][21] ), .S0(n9196), .S1(n9197), .Q(n6780) );
  MUX41X1 U4783 ( .IN1(\R[3][19] ), .IN3(\R[1][19] ), .IN2(\R[2][19] ), .IN4(
        \R[0][19] ), .S0(n9196), .S1(n9197), .Q(n6776) );
  MUX41X1 U4784 ( .IN1(\R[3][17] ), .IN3(\R[1][17] ), .IN2(\R[2][17] ), .IN4(
        \R[0][17] ), .S0(n9196), .S1(n9197), .Q(n6772) );
  MUX41X1 U4785 ( .IN1(\R[3][15] ), .IN3(\R[1][15] ), .IN2(\R[2][15] ), .IN4(
        \R[0][15] ), .S0(n9196), .S1(n9197), .Q(n6768) );
  INVX0 U4786 ( .INP(n9197), .ZN(n6801) );
  INVX0 U4787 ( .INP(n9197), .ZN(n6802) );
  INVX0 U4788 ( .INP(n9197), .ZN(n6803) );
  INVX0 U4789 ( .INP(n9197), .ZN(n6804) );
  INVX0 U4790 ( .INP(n9197), .ZN(n6805) );
  INVX0 U4791 ( .INP(n9197), .ZN(n6806) );
  INVX0 U4792 ( .INP(n9197), .ZN(n6807) );
  MUX41X1 U4793 ( .IN1(\R[3][1] ), .IN3(\R[1][1] ), .IN2(\R[2][1] ), .IN4(
        \R[0][1] ), .S0(n9193), .S1(n9194), .Q(n6811) );
  MUX41X1 U4794 ( .IN1(\R[3][3] ), .IN3(\R[1][3] ), .IN2(\R[2][3] ), .IN4(
        \R[0][3] ), .S0(n9193), .S1(n9194), .Q(n6815) );
  MUX41X1 U4795 ( .IN1(\R[3][5] ), .IN3(\R[1][5] ), .IN2(\R[2][5] ), .IN4(
        \R[0][5] ), .S0(n9193), .S1(n9194), .Q(n6819) );
  MUX41X1 U4796 ( .IN1(\R[3][8] ), .IN3(\R[1][8] ), .IN2(\R[2][8] ), .IN4(
        \R[0][8] ), .S0(n9193), .S1(n9194), .Q(n6825) );
  MUX41X1 U4797 ( .IN1(\R[3][10] ), .IN3(\R[1][10] ), .IN2(\R[2][10] ), .IN4(
        \R[0][10] ), .S0(n9193), .S1(n9194), .Q(n6829) );
  INVX0 U4798 ( .INP(n9194), .ZN(n6877) );
  MUX41X1 U4799 ( .IN1(\R[3][12] ), .IN3(\R[1][12] ), .IN2(\R[2][12] ), .IN4(
        \R[0][12] ), .S0(n9193), .S1(n9194), .Q(n6833) );
  INVX0 U4800 ( .INP(n9194), .ZN(n6876) );
  MUX41X1 U4801 ( .IN1(\R[3][14] ), .IN3(\R[1][14] ), .IN2(\R[2][14] ), .IN4(
        \R[0][14] ), .S0(n9193), .S1(n9194), .Q(n6837) );
  INVX0 U4802 ( .INP(n9194), .ZN(n6875) );
  MUX41X1 U4803 ( .IN1(\R[3][16] ), .IN3(\R[1][16] ), .IN2(\R[2][16] ), .IN4(
        \R[0][16] ), .S0(n9193), .S1(n9194), .Q(n6841) );
  INVX0 U4804 ( .INP(n9194), .ZN(n6874) );
  INVX0 U4805 ( .INP(n9194), .ZN(n6873) );
  INVX0 U4806 ( .INP(n9194), .ZN(n6872) );
  OA21X1 U4807 ( .IN1(N1865), .IN2(n5753), .IN3(n6039), .Q(n6038) );
  OA21X1 U4808 ( .IN1(N1867), .IN2(n5753), .IN3(n5983), .Q(n5982) );
  OA21X1 U4809 ( .IN1(N1869), .IN2(n5753), .IN3(n5927), .Q(n5926) );
  OA21X1 U4810 ( .IN1(N1874), .IN2(n5753), .IN3(n6347), .Q(n6346) );
  OA21X1 U4811 ( .IN1(N1875), .IN2(n5753), .IN3(n6319), .Q(n6318) );
  OA21X1 U4812 ( .IN1(N1876), .IN2(n5753), .IN3(n6095), .Q(n6094) );
  OA21X1 U4813 ( .IN1(N1877), .IN2(n5753), .IN3(n6291), .Q(n6290) );
  OA21X1 U4814 ( .IN1(N1879), .IN2(n5753), .IN3(n6235), .Q(n6234) );
  OA21X1 U4815 ( .IN1(N1880), .IN2(n5753), .IN3(n6207), .Q(n6206) );
  OA21X1 U4816 ( .IN1(N1881), .IN2(n5753), .IN3(n6179), .Q(n6178) );
  OA21X1 U4817 ( .IN1(N1882), .IN2(n5753), .IN3(n6151), .Q(n6150) );
  OA21X1 U4818 ( .IN1(N1883), .IN2(n5753), .IN3(n6123), .Q(n6122) );
  OA21X1 U4819 ( .IN1(N1885), .IN2(n5753), .IN3(n6401), .Q(n6400) );
  OA21X1 U4820 ( .IN1(N1886), .IN2(n5753), .IN3(n6374), .Q(n6373) );
  OA21X1 U4821 ( .IN1(N1887), .IN2(n5753), .IN3(n6457), .Q(n6456) );
  OA21X1 U4822 ( .IN1(N1892), .IN2(n5753), .IN3(n6536), .Q(n6535) );
  OA21X1 U4823 ( .IN1(N1893), .IN2(n5753), .IN3(n6510), .Q(n6509) );
  OA21X1 U4824 ( .IN1(N1894), .IN2(n5753), .IN3(n6484), .Q(n6483) );
  INVX0 U4825 ( .INP(n3700), .ZN(n7015) );
  INVX0 U4826 ( .INP(n3700), .ZN(n7016) );
  INVX0 U4827 ( .INP(n3700), .ZN(n7017) );
  INVX0 U4828 ( .INP(n3700), .ZN(n7018) );
  INVX0 U4829 ( .INP(n3700), .ZN(n7019) );
  INVX0 U4830 ( .INP(n3700), .ZN(n7020) );
  INVX0 U4831 ( .INP(n3700), .ZN(n7021) );
  INVX0 U4832 ( .INP(n3700), .ZN(n7022) );
  INVX0 U4833 ( .INP(n3700), .ZN(n7023) );
  INVX0 U4834 ( .INP(n3700), .ZN(n7024) );
  INVX0 U4835 ( .INP(n3700), .ZN(n7025) );
  INVX0 U4836 ( .INP(n3700), .ZN(n7026) );
  OA21X1 U4837 ( .IN1(N1864), .IN2(n5696), .IN3(n6067), .Q(n6066) );
  OA21X1 U4838 ( .IN1(N1866), .IN2(n5696), .IN3(n6011), .Q(n6010) );
  OA21X1 U4839 ( .IN1(N1868), .IN2(n5696), .IN3(n5955), .Q(n5954) );
  OA21X1 U4840 ( .IN1(N1870), .IN2(n5696), .IN3(n5899), .Q(n5898) );
  OA21X1 U4841 ( .IN1(N1871), .IN2(n5696), .IN3(n5871), .Q(n5870) );
  OA21X1 U4842 ( .IN1(N1872), .IN2(n5696), .IN3(n5843), .Q(n5842) );
  OA21X1 U4843 ( .IN1(N1873), .IN2(n5696), .IN3(n5815), .Q(n5814) );
  OA21X1 U4844 ( .IN1(N1878), .IN2(n5696), .IN3(n6263), .Q(n6262) );
  OA21X1 U4845 ( .IN1(N1884), .IN2(n5696), .IN3(n6429), .Q(n6428) );
  OA21X1 U4846 ( .IN1(N1888), .IN2(n5696), .IN3(n6640), .Q(n6639) );
  OA21X1 U4847 ( .IN1(N1889), .IN2(n5696), .IN3(n6614), .Q(n6613) );
  OA21X1 U4848 ( .IN1(N1890), .IN2(n5696), .IN3(n6588), .Q(n6587) );
  OA21X1 U4849 ( .IN1(N1891), .IN2(n5696), .IN3(n6562), .Q(n6561) );
  OA21X1 U4850 ( .IN1(N1895), .IN2(n5696), .IN3(n6665), .Q(n6664) );
  INVX0 U4851 ( .INP(n3723), .ZN(n5724) );
  INVX0 U4852 ( .INP(n3723), .ZN(n5725) );
  INVX0 U4853 ( .INP(n3723), .ZN(n5726) );
  INVX0 U4854 ( .INP(n3723), .ZN(n5727) );
  INVX0 U4855 ( .INP(n3723), .ZN(n5728) );
  INVX0 U4856 ( .INP(n3723), .ZN(n5729) );
  INVX0 U4857 ( .INP(n3723), .ZN(n5730) );
  INVX0 U4858 ( .INP(n3723), .ZN(n5731) );
  INVX0 U4859 ( .INP(n3723), .ZN(n5732) );
  INVX0 U4860 ( .INP(n3723), .ZN(n5733) );
  INVX0 U4861 ( .INP(n3723), .ZN(n5734) );
  INVX0 U4862 ( .INP(n3723), .ZN(n5735) );
  INVX0 U4863 ( .INP(n3723), .ZN(n5736) );
  INVX0 U4864 ( .INP(n3723), .ZN(n5737) );
  INVX0 U4865 ( .INP(n3723), .ZN(n5738) );
  INVX0 U4866 ( .INP(n3723), .ZN(n5739) );
  INVX0 U4867 ( .INP(n3723), .ZN(n5740) );
  INVX0 U4868 ( .INP(n3723), .ZN(n5741) );
  INVX0 U4869 ( .INP(n3723), .ZN(n5742) );
  INVX0 U4870 ( .INP(n3723), .ZN(n5743) );
  INVX0 U4871 ( .INP(n3723), .ZN(n5744) );
  INVX0 U4872 ( .INP(n3721), .ZN(n5745) );
  INVX0 U4873 ( .INP(n3721), .ZN(n5746) );
  INVX0 U4874 ( .INP(n3721), .ZN(n5747) );
  INVX0 U4875 ( .INP(n3721), .ZN(n5748) );
  INVX0 U4876 ( .INP(n3721), .ZN(n5749) );
  INVX0 U4877 ( .INP(n3721), .ZN(n5750) );
  INVX0 U4878 ( .INP(n3721), .ZN(n5751) );
  INVX0 U4879 ( .INP(n3721), .ZN(n5752) );
  INVX0 U4880 ( .INP(n3721), .ZN(n5753) );
  INVX0 U4881 ( .INP(n5784), .ZN(n5754) );
  INVX0 U4882 ( .INP(n5783), .ZN(n5755) );
  INVX0 U4883 ( .INP(n5784), .ZN(n5756) );
  INVX0 U4884 ( .INP(n5784), .ZN(n5757) );
  INVX0 U4885 ( .INP(n5784), .ZN(n5758) );
  INVX0 U4886 ( .INP(n5783), .ZN(n5759) );
  INVX0 U4887 ( .INP(n5783), .ZN(n5760) );
  INVX0 U4888 ( .INP(n5783), .ZN(n5761) );
  INVX0 U4889 ( .INP(n5782), .ZN(n5762) );
  INVX0 U4890 ( .INP(n5782), .ZN(n5763) );
  INVX0 U4891 ( .INP(n5782), .ZN(n5764) );
  INVX0 U4892 ( .INP(n5782), .ZN(n5765) );
  INVX0 U4893 ( .INP(n5781), .ZN(n5766) );
  INVX0 U4894 ( .INP(n5780), .ZN(n5767) );
  INVX0 U4895 ( .INP(n5781), .ZN(n5768) );
  INVX0 U4896 ( .INP(n5781), .ZN(n5769) );
  INVX0 U4897 ( .INP(n5781), .ZN(n5770) );
  INVX0 U4898 ( .INP(n5780), .ZN(n5771) );
  INVX0 U4899 ( .INP(n5780), .ZN(n5772) );
  INVX0 U4900 ( .INP(n5780), .ZN(n5773) );
  INVX0 U4901 ( .INP(n5786), .ZN(n5774) );
  INVX0 U4902 ( .INP(n5785), .ZN(n5775) );
  INVX0 U4903 ( .INP(n5784), .ZN(n5776) );
  INVX0 U4904 ( .INP(n5780), .ZN(n5777) );
  INVX0 U4905 ( .INP(n5786), .ZN(n5778) );
  INVX0 U4906 ( .INP(n5785), .ZN(n5779) );
  INVX0 U4907 ( .INP(\U3/U85/Z_4 ), .ZN(n5780) );
  INVX0 U4908 ( .INP(\U3/U85/Z_4 ), .ZN(n5781) );
  INVX0 U4909 ( .INP(\U3/U85/Z_4 ), .ZN(n5782) );
  INVX0 U4910 ( .INP(\U3/U85/Z_4 ), .ZN(n5783) );
  INVX0 U4911 ( .INP(\U3/U85/Z_4 ), .ZN(n5784) );
  INVX0 U4912 ( .INP(\U3/U85/Z_4 ), .ZN(n5785) );
  INVX0 U4913 ( .INP(\U3/U85/Z_4 ), .ZN(n5786) );
  MUX21X1 U4914 ( .IN1(N4799), .IN2(N4868), .S(n5757), .Q(n5797) );
  MUX21X1 U4915 ( .IN1(N1757), .IN2(n5797), .S(n5736), .Q(n5798) );
  MUX21X1 U4916 ( .IN1(N4601), .IN2(N1757), .S(n5768), .Q(n5799) );
  MUX21X1 U4917 ( .IN1(n516), .IN2(N1757), .S(n5766), .Q(n5800) );
  MUX21X1 U4918 ( .IN1(N4360), .IN2(ID_imm_offset[10]), .S(n5766), .Q(n5801)
         );
  MUX41X1 U4919 ( .IN1(n5801), .IN3(N5282), .IN2(n5800), .IN4(n5799), .S0(
        n5750), .S1(n5724), .Q(n5802) );
  MUX21X1 U4920 ( .IN1(n5802), .IN2(n5798), .S(n5787), .Q(n5803) );
  MUX21X1 U4921 ( .IN1(N4733), .IN2(N4766), .S(n5736), .Q(n5804) );
  MUX21X1 U4922 ( .IN1(n5804), .IN2(N1757), .S(n5767), .Q(n5805) );
  MUX21X1 U4923 ( .IN1(n516), .IN2(N5217), .S(n5736), .Q(n5806) );
  MUX21X1 U4924 ( .IN1(N3007), .IN2(N4132), .S(n5767), .Q(n5807) );
  MUX21X1 U4925 ( .IN1(n5807), .IN2(n5723), .S(n5736), .Q(n5808) );
  MUX41X1 U4926 ( .IN1(n5808), .IN3(n5805), .IN2(n5806), .IN4(n4433), .S0(
        n5792), .S1(n5745), .Q(n5809) );
  MUX21X1 U4927 ( .IN1(N1757), .IN2(n516), .S(n5767), .Q(n5810) );
  MUX21X1 U4928 ( .IN1(N4503), .IN2(N4536), .S(n5767), .Q(n5811) );
  MUX21X1 U4929 ( .IN1(N1790), .IN2(N1822), .S(n5767), .Q(n5812) );
  MUX41X1 U4930 ( .IN1(n5799), .IN3(n5810), .IN2(n5812), .IN4(n5811), .S0(
        n5750), .S1(n5724), .Q(n5813) );
  MUX21X1 U4931 ( .IN1(n5814), .IN2(n5813), .S(n5787), .Q(n5816) );
  MUX41X1 U4932 ( .IN1(N1822), .IN3(N1757), .IN2(N4733), .IN4(N4766), .S0(
        n5744), .S1(n5754), .Q(n5817) );
  MUX21X1 U4933 ( .IN1(n5811), .IN2(N4556), .S(n5736), .Q(n5818) );
  MUX21X1 U4934 ( .IN1(N4902), .IN2(N4970), .S(n5767), .Q(n5819) );
  AND2X1 U4935 ( .IN1(N5003), .IN2(n5779), .Q(n5820) );
  MUX21X1 U4936 ( .IN1(n5819), .IN2(n5820), .S(n5736), .Q(n5821) );
  MUX21X1 U4937 ( .IN1(n516), .IN2(N1757), .S(n5736), .Q(n5822) );
  MUX21X1 U4938 ( .IN1(n403), .IN2(n5822), .S(n5767), .Q(n5823) );
  MUX41X1 U4939 ( .IN1(n5823), .IN3(n5818), .IN2(n5821), .IN4(n5817), .S0(
        n5796), .S1(n5745), .Q(n5824) );
  MUX41X1 U4940 ( .IN1(n5824), .IN3(n5816), .IN2(n5809), .IN4(n5803), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5644) );
  MUX21X1 U4941 ( .IN1(N4800), .IN2(N4869), .S(n5767), .Q(n5825) );
  MUX21X1 U4942 ( .IN1(N1758), .IN2(n5825), .S(n5736), .Q(n5826) );
  MUX21X1 U4943 ( .IN1(N4602), .IN2(N1758), .S(n5767), .Q(n5827) );
  MUX21X1 U4944 ( .IN1(n515), .IN2(N1758), .S(n5767), .Q(n5828) );
  MUX21X1 U4945 ( .IN1(N4359), .IN2(ID_imm_offset[10]), .S(n5767), .Q(n5829)
         );
  MUX41X1 U4946 ( .IN1(n5829), .IN3(N5283), .IN2(n5828), .IN4(n5827), .S0(
        n5750), .S1(n5724), .Q(n5830) );
  MUX21X1 U4947 ( .IN1(n5830), .IN2(n5826), .S(n5787), .Q(n5831) );
  MUX21X1 U4948 ( .IN1(N4734), .IN2(N4767), .S(n5736), .Q(n5832) );
  MUX21X1 U4949 ( .IN1(n5832), .IN2(N1758), .S(n5767), .Q(n5833) );
  MUX21X1 U4950 ( .IN1(n515), .IN2(N5218), .S(n5735), .Q(n5834) );
  MUX21X1 U4951 ( .IN1(N3008), .IN2(N4133), .S(n5767), .Q(n5835) );
  MUX21X1 U4952 ( .IN1(n5835), .IN2(n5723), .S(n5735), .Q(n5836) );
  MUX41X1 U4953 ( .IN1(n5836), .IN3(n5833), .IN2(n5834), .IN4(n4432), .S0(
        n5796), .S1(n5745), .Q(n5837) );
  MUX21X1 U4954 ( .IN1(N1758), .IN2(n515), .S(n5767), .Q(n5838) );
  MUX21X1 U4955 ( .IN1(N4504), .IN2(N4537), .S(n5767), .Q(n5839) );
  MUX21X1 U4956 ( .IN1(N1791), .IN2(N1823), .S(n5767), .Q(n5840) );
  MUX41X1 U4957 ( .IN1(n5827), .IN3(n5838), .IN2(n5840), .IN4(n5839), .S0(
        n5750), .S1(n5724), .Q(n5841) );
  MUX21X1 U4958 ( .IN1(n5842), .IN2(n5841), .S(n5787), .Q(n5844) );
  MUX41X1 U4959 ( .IN1(N1823), .IN3(N1758), .IN2(N4734), .IN4(N4767), .S0(
        n5744), .S1(n5754), .Q(n5845) );
  MUX21X1 U4960 ( .IN1(n5839), .IN2(N4555), .S(n5735), .Q(n5846) );
  MUX21X1 U4961 ( .IN1(N4903), .IN2(N4971), .S(n5767), .Q(n5847) );
  AND2X1 U4962 ( .IN1(N5004), .IN2(n5778), .Q(n5848) );
  MUX21X1 U4963 ( .IN1(n5847), .IN2(n5848), .S(n5735), .Q(n5849) );
  MUX21X1 U4964 ( .IN1(n515), .IN2(N1758), .S(n5735), .Q(n5850) );
  MUX21X1 U4965 ( .IN1(n402), .IN2(n5850), .S(n5767), .Q(n5851) );
  MUX41X1 U4966 ( .IN1(n5851), .IN3(n5846), .IN2(n5849), .IN4(n5845), .S0(
        n5796), .S1(n5745), .Q(n5852) );
  MUX41X1 U4967 ( .IN1(n5852), .IN3(n5844), .IN2(n5837), .IN4(n5831), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5645) );
  MUX21X1 U4968 ( .IN1(N4801), .IN2(N4870), .S(n5768), .Q(n5853) );
  MUX21X1 U4969 ( .IN1(N1759), .IN2(n5853), .S(n5735), .Q(n5854) );
  MUX21X1 U4970 ( .IN1(N4603), .IN2(N1759), .S(n5768), .Q(n5855) );
  MUX21X1 U4971 ( .IN1(n514), .IN2(N1759), .S(n5768), .Q(n5856) );
  MUX21X1 U4972 ( .IN1(N4358), .IN2(ID_imm_offset[10]), .S(n5768), .Q(n5857)
         );
  MUX41X1 U4973 ( .IN1(n5857), .IN3(N5284), .IN2(n5856), .IN4(n5855), .S0(
        n5750), .S1(n5725), .Q(n5858) );
  MUX21X1 U4974 ( .IN1(n5858), .IN2(n5854), .S(n5787), .Q(n5859) );
  MUX21X1 U4975 ( .IN1(N4735), .IN2(N4768), .S(n5735), .Q(n5860) );
  MUX21X1 U4976 ( .IN1(n5860), .IN2(N1759), .S(n5768), .Q(n5861) );
  MUX21X1 U4977 ( .IN1(n514), .IN2(N5219), .S(n5735), .Q(n5862) );
  MUX21X1 U4978 ( .IN1(N3009), .IN2(N4134), .S(n5768), .Q(n5863) );
  MUX21X1 U4979 ( .IN1(n5863), .IN2(n5723), .S(n5735), .Q(n5864) );
  MUX41X1 U4980 ( .IN1(n5864), .IN3(n5861), .IN2(n5862), .IN4(n4431), .S0(
        n5796), .S1(n5745), .Q(n5865) );
  MUX21X1 U4981 ( .IN1(N1759), .IN2(n514), .S(n5768), .Q(n5866) );
  MUX21X1 U4982 ( .IN1(N4505), .IN2(N4538), .S(n5772), .Q(n5867) );
  MUX21X1 U4983 ( .IN1(N1792), .IN2(N1824), .S(n5768), .Q(n5868) );
  MUX41X1 U4984 ( .IN1(n5855), .IN3(n5866), .IN2(n5868), .IN4(n5867), .S0(
        n5750), .S1(n5725), .Q(n5869) );
  MUX21X1 U4985 ( .IN1(n5870), .IN2(n5869), .S(n5787), .Q(n5872) );
  MUX41X1 U4986 ( .IN1(N1824), .IN3(N1759), .IN2(N4735), .IN4(N4768), .S0(
        n5744), .S1(n5756), .Q(n5873) );
  MUX21X1 U4987 ( .IN1(n5867), .IN2(N4554), .S(n5735), .Q(n5874) );
  MUX21X1 U4988 ( .IN1(N4904), .IN2(N4972), .S(n5768), .Q(n5875) );
  AND2X1 U4989 ( .IN1(N5005), .IN2(n5778), .Q(n5876) );
  MUX21X1 U4990 ( .IN1(n5875), .IN2(n5876), .S(n5735), .Q(n5877) );
  MUX21X1 U4991 ( .IN1(n514), .IN2(N1759), .S(n5735), .Q(n5878) );
  MUX21X1 U4992 ( .IN1(n401), .IN2(n5878), .S(n5768), .Q(n5879) );
  MUX41X1 U4993 ( .IN1(n5879), .IN3(n5874), .IN2(n5877), .IN4(n5873), .S0(
        n5796), .S1(n5746), .Q(n5880) );
  MUX41X1 U4994 ( .IN1(n5880), .IN3(n5872), .IN2(n5865), .IN4(n5859), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5646) );
  MUX21X1 U4995 ( .IN1(N4802), .IN2(N4871), .S(n5768), .Q(n5881) );
  MUX21X1 U4996 ( .IN1(N1760), .IN2(n5881), .S(n5735), .Q(n5882) );
  MUX21X1 U4997 ( .IN1(N4604), .IN2(N1760), .S(n5768), .Q(n5883) );
  MUX21X1 U4998 ( .IN1(n513), .IN2(N1760), .S(n5768), .Q(n5884) );
  MUX21X1 U4999 ( .IN1(N4357), .IN2(ID_imm_offset[10]), .S(n5768), .Q(n5885)
         );
  MUX41X1 U5000 ( .IN1(n5885), .IN3(N5285), .IN2(n5884), .IN4(n5883), .S0(
        n5751), .S1(n5725), .Q(n5886) );
  MUX21X1 U5001 ( .IN1(n5886), .IN2(n5882), .S(n5787), .Q(n5887) );
  MUX21X1 U5002 ( .IN1(N4736), .IN2(N4769), .S(n5735), .Q(n5888) );
  MUX21X1 U5003 ( .IN1(n5888), .IN2(N1760), .S(n5768), .Q(n5889) );
  MUX21X1 U5004 ( .IN1(n513), .IN2(N5220), .S(n5735), .Q(n5890) );
  MUX21X1 U5005 ( .IN1(N3010), .IN2(N4135), .S(n5768), .Q(n5891) );
  MUX21X1 U5006 ( .IN1(n5891), .IN2(n5723), .S(n5735), .Q(n5892) );
  MUX41X1 U5007 ( .IN1(n5892), .IN3(n5889), .IN2(n5890), .IN4(n4430), .S0(
        n5796), .S1(n5746), .Q(n5893) );
  MUX21X1 U5008 ( .IN1(N1760), .IN2(n513), .S(n5768), .Q(n5894) );
  MUX21X1 U5009 ( .IN1(N4506), .IN2(N4539), .S(n5769), .Q(n5895) );
  MUX21X1 U5010 ( .IN1(N1793), .IN2(N1825), .S(n5769), .Q(n5896) );
  MUX41X1 U5011 ( .IN1(n5883), .IN3(n5894), .IN2(n5896), .IN4(n5895), .S0(
        n5751), .S1(n5726), .Q(n5897) );
  MUX21X1 U5012 ( .IN1(n5898), .IN2(n5897), .S(n5787), .Q(n5900) );
  MUX41X1 U5013 ( .IN1(N1825), .IN3(N1760), .IN2(N4736), .IN4(N4769), .S0(
        n5744), .S1(n5755), .Q(n5901) );
  MUX21X1 U5014 ( .IN1(n5895), .IN2(N4553), .S(n5735), .Q(n5902) );
  MUX21X1 U5015 ( .IN1(N4905), .IN2(N4973), .S(n5769), .Q(n5903) );
  AND2X1 U5016 ( .IN1(N5006), .IN2(n5779), .Q(n5904) );
  MUX21X1 U5017 ( .IN1(n5903), .IN2(n5904), .S(n5735), .Q(n5905) );
  MUX21X1 U5018 ( .IN1(n513), .IN2(N1760), .S(n5734), .Q(n5906) );
  MUX21X1 U5019 ( .IN1(n400), .IN2(n5906), .S(n5769), .Q(n5907) );
  MUX41X1 U5020 ( .IN1(n5907), .IN3(n5902), .IN2(n5905), .IN4(n5901), .S0(
        n5796), .S1(n5746), .Q(n5908) );
  MUX41X1 U5021 ( .IN1(n5908), .IN3(n5900), .IN2(n5893), .IN4(n5887), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5647) );
  MUX21X1 U5022 ( .IN1(N4803), .IN2(N4872), .S(n5769), .Q(n5909) );
  MUX21X1 U5023 ( .IN1(N1761), .IN2(n5909), .S(n5734), .Q(n5910) );
  MUX21X1 U5024 ( .IN1(N4605), .IN2(N1761), .S(n5769), .Q(n5911) );
  MUX21X1 U5025 ( .IN1(n512), .IN2(N1761), .S(n5769), .Q(n5912) );
  MUX21X1 U5026 ( .IN1(N4356), .IN2(ID_imm_offset[10]), .S(n5769), .Q(n5913)
         );
  MUX41X1 U5027 ( .IN1(n5913), .IN3(N5286), .IN2(n5912), .IN4(n5911), .S0(
        n5751), .S1(n5727), .Q(n5914) );
  MUX21X1 U5028 ( .IN1(n5914), .IN2(n5910), .S(n5788), .Q(n5915) );
  MUX21X1 U5029 ( .IN1(N4737), .IN2(N4770), .S(n5734), .Q(n5916) );
  MUX21X1 U5030 ( .IN1(n5916), .IN2(N1761), .S(n5769), .Q(n5917) );
  MUX21X1 U5031 ( .IN1(n512), .IN2(N5221), .S(n5734), .Q(n5918) );
  MUX21X1 U5032 ( .IN1(N3011), .IN2(N4136), .S(n5769), .Q(n5919) );
  MUX21X1 U5033 ( .IN1(n5919), .IN2(n5723), .S(n5734), .Q(n5920) );
  MUX41X1 U5034 ( .IN1(n5920), .IN3(n5917), .IN2(n5918), .IN4(n4429), .S0(
        n5796), .S1(n5746), .Q(n5921) );
  MUX21X1 U5035 ( .IN1(N1761), .IN2(n512), .S(n5769), .Q(n5922) );
  MUX21X1 U5036 ( .IN1(N4507), .IN2(N4540), .S(n5769), .Q(n5923) );
  MUX21X1 U5037 ( .IN1(N1794), .IN2(N1826), .S(n5769), .Q(n5924) );
  MUX41X1 U5038 ( .IN1(n5911), .IN3(n5922), .IN2(n5924), .IN4(n5923), .S0(
        n5750), .S1(n5727), .Q(n5925) );
  MUX21X1 U5039 ( .IN1(n5926), .IN2(n5925), .S(n5788), .Q(n5928) );
  MUX41X1 U5040 ( .IN1(N1826), .IN3(N1761), .IN2(N4737), .IN4(N4770), .S0(
        n5695), .S1(n5756), .Q(n5929) );
  MUX21X1 U5041 ( .IN1(n5923), .IN2(N4552), .S(n5734), .Q(n5930) );
  MUX21X1 U5042 ( .IN1(N4906), .IN2(N4974), .S(n5769), .Q(n5931) );
  AND2X1 U5043 ( .IN1(N5007), .IN2(n5779), .Q(n5932) );
  MUX21X1 U5044 ( .IN1(n5931), .IN2(n5932), .S(n5734), .Q(n5933) );
  MUX21X1 U5045 ( .IN1(n512), .IN2(N1761), .S(n5734), .Q(n5934) );
  MUX21X1 U5046 ( .IN1(n399), .IN2(n5934), .S(n5769), .Q(n5935) );
  MUX41X1 U5047 ( .IN1(n5935), .IN3(n5930), .IN2(n5933), .IN4(n5929), .S0(
        n5796), .S1(n5747), .Q(n5936) );
  MUX41X1 U5048 ( .IN1(n5936), .IN3(n5928), .IN2(n5921), .IN4(n5915), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5648) );
  MUX21X1 U5049 ( .IN1(N4804), .IN2(N4873), .S(n5769), .Q(n5937) );
  MUX21X1 U5050 ( .IN1(N1762), .IN2(n5937), .S(n5734), .Q(n5938) );
  MUX21X1 U5051 ( .IN1(N4606), .IN2(N1762), .S(n5769), .Q(n5939) );
  MUX21X1 U5052 ( .IN1(n511), .IN2(N1762), .S(n5769), .Q(n5940) );
  MUX21X1 U5053 ( .IN1(N4355), .IN2(ID_imm_offset[10]), .S(n5770), .Q(n5941)
         );
  MUX41X1 U5054 ( .IN1(n5941), .IN3(N5287), .IN2(n5940), .IN4(n5939), .S0(
        n5751), .S1(n5728), .Q(n5942) );
  MUX21X1 U5055 ( .IN1(n5942), .IN2(n5938), .S(n5788), .Q(n5943) );
  MUX21X1 U5056 ( .IN1(N4738), .IN2(N4771), .S(n5734), .Q(n5944) );
  MUX21X1 U5057 ( .IN1(n5944), .IN2(N1762), .S(n5770), .Q(n5945) );
  MUX21X1 U5058 ( .IN1(n511), .IN2(N5222), .S(n5734), .Q(n5946) );
  MUX21X1 U5059 ( .IN1(N3012), .IN2(N4137), .S(n5770), .Q(n5947) );
  MUX21X1 U5060 ( .IN1(n5947), .IN2(n5723), .S(n5734), .Q(n5948) );
  MUX41X1 U5061 ( .IN1(n5948), .IN3(n5945), .IN2(n5946), .IN4(n4428), .S0(
        n5795), .S1(n5746), .Q(n5949) );
  MUX21X1 U5062 ( .IN1(N1762), .IN2(n511), .S(n5770), .Q(n5950) );
  MUX21X1 U5063 ( .IN1(N4508), .IN2(N4541), .S(n5770), .Q(n5951) );
  MUX21X1 U5064 ( .IN1(N1795), .IN2(N1827), .S(n5770), .Q(n5952) );
  MUX41X1 U5065 ( .IN1(n5939), .IN3(n5950), .IN2(n5952), .IN4(n5951), .S0(
        n5750), .S1(n5728), .Q(n5953) );
  MUX21X1 U5066 ( .IN1(n5954), .IN2(n5953), .S(n5788), .Q(n5956) );
  MUX41X1 U5067 ( .IN1(N1827), .IN3(N1762), .IN2(N4738), .IN4(N4771), .S0(
        n5743), .S1(n5756), .Q(n5957) );
  MUX21X1 U5068 ( .IN1(n5951), .IN2(N4551), .S(n5734), .Q(n5958) );
  MUX21X1 U5069 ( .IN1(N4907), .IN2(N4975), .S(n5770), .Q(n5959) );
  AND2X1 U5070 ( .IN1(N5008), .IN2(n5778), .Q(n5960) );
  MUX21X1 U5071 ( .IN1(n5959), .IN2(n5960), .S(n5734), .Q(n5961) );
  MUX21X1 U5072 ( .IN1(n511), .IN2(N1762), .S(n5734), .Q(n5962) );
  MUX21X1 U5073 ( .IN1(n398), .IN2(n5962), .S(n5770), .Q(n5963) );
  MUX41X1 U5074 ( .IN1(n5963), .IN3(n5958), .IN2(n5961), .IN4(n5957), .S0(
        n5795), .S1(n5747), .Q(n5964) );
  MUX41X1 U5075 ( .IN1(n5964), .IN3(n5956), .IN2(n5949), .IN4(n5943), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5649) );
  MUX21X1 U5076 ( .IN1(N4805), .IN2(N4874), .S(n5770), .Q(n5965) );
  MUX21X1 U5077 ( .IN1(N1763), .IN2(n5965), .S(n5734), .Q(n5966) );
  MUX21X1 U5078 ( .IN1(N4607), .IN2(N1763), .S(n5770), .Q(n5967) );
  MUX21X1 U5079 ( .IN1(n510), .IN2(N1763), .S(n5770), .Q(n5968) );
  MUX21X1 U5080 ( .IN1(N4354), .IN2(ID_imm_offset[10]), .S(n5770), .Q(n5969)
         );
  MUX41X1 U5081 ( .IN1(n5969), .IN3(N5288), .IN2(n5968), .IN4(n5967), .S0(
        n5750), .S1(n5727), .Q(n5970) );
  MUX21X1 U5082 ( .IN1(n5970), .IN2(n5966), .S(n5788), .Q(n5971) );
  MUX21X1 U5083 ( .IN1(N4739), .IN2(N4772), .S(n5734), .Q(n5972) );
  MUX21X1 U5084 ( .IN1(n5972), .IN2(N1763), .S(n5770), .Q(n5973) );
  MUX21X1 U5085 ( .IN1(n510), .IN2(N5223), .S(n5734), .Q(n5974) );
  MUX21X1 U5086 ( .IN1(N3013), .IN2(N4138), .S(n5770), .Q(n5975) );
  MUX21X1 U5087 ( .IN1(n5975), .IN2(n5723), .S(n5733), .Q(n5976) );
  MUX41X1 U5088 ( .IN1(n5976), .IN3(n5973), .IN2(n5974), .IN4(n4427), .S0(
        n5795), .S1(n5747), .Q(n5977) );
  MUX21X1 U5089 ( .IN1(N1763), .IN2(n510), .S(n5770), .Q(n5978) );
  MUX21X1 U5090 ( .IN1(N4509), .IN2(N4542), .S(n5770), .Q(n5979) );
  MUX21X1 U5091 ( .IN1(N1796), .IN2(N1828), .S(n5770), .Q(n5980) );
  MUX41X1 U5092 ( .IN1(n5967), .IN3(n5978), .IN2(n5980), .IN4(n5979), .S0(
        n5751), .S1(n5728), .Q(n5981) );
  MUX21X1 U5093 ( .IN1(n5982), .IN2(n5981), .S(n5788), .Q(n5984) );
  MUX41X1 U5094 ( .IN1(N1828), .IN3(N1763), .IN2(N4739), .IN4(N4772), .S0(
        n5744), .S1(n5756), .Q(n5985) );
  MUX21X1 U5095 ( .IN1(n5979), .IN2(N4550), .S(n5733), .Q(n5986) );
  MUX21X1 U5096 ( .IN1(N4908), .IN2(N4976), .S(n5770), .Q(n5987) );
  AND2X1 U5097 ( .IN1(N5009), .IN2(n5778), .Q(n5988) );
  MUX21X1 U5098 ( .IN1(n5987), .IN2(n5988), .S(n5733), .Q(n5989) );
  MUX21X1 U5099 ( .IN1(n510), .IN2(N1763), .S(n5733), .Q(n5990) );
  MUX21X1 U5100 ( .IN1(n397), .IN2(n5990), .S(n5771), .Q(n5991) );
  MUX41X1 U5101 ( .IN1(n5991), .IN3(n5986), .IN2(n5989), .IN4(n5985), .S0(
        n5795), .S1(n5747), .Q(n5992) );
  MUX41X1 U5102 ( .IN1(n5992), .IN3(n5984), .IN2(n5977), .IN4(n5971), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5650) );
  MUX21X1 U5103 ( .IN1(N4806), .IN2(N4875), .S(n5771), .Q(n5993) );
  MUX21X1 U5104 ( .IN1(N1764), .IN2(n5993), .S(n5733), .Q(n5994) );
  MUX21X1 U5105 ( .IN1(N4608), .IN2(N1764), .S(n5771), .Q(n5995) );
  MUX21X1 U5106 ( .IN1(n509), .IN2(N1764), .S(n5771), .Q(n5996) );
  MUX21X1 U5107 ( .IN1(N4353), .IN2(ID_imm_offset[10]), .S(n5771), .Q(n5997)
         );
  MUX41X1 U5108 ( .IN1(n5997), .IN3(N5289), .IN2(n5996), .IN4(n5995), .S0(
        n5750), .S1(n5729), .Q(n5998) );
  MUX21X1 U5109 ( .IN1(n5998), .IN2(n5994), .S(n5788), .Q(n5999) );
  MUX21X1 U5110 ( .IN1(N4740), .IN2(N4773), .S(n5733), .Q(n6000) );
  MUX21X1 U5111 ( .IN1(n6000), .IN2(N1764), .S(n5771), .Q(n6001) );
  MUX21X1 U5112 ( .IN1(n509), .IN2(N5224), .S(n5733), .Q(n6002) );
  MUX21X1 U5113 ( .IN1(N3014), .IN2(N4139), .S(n5771), .Q(n6003) );
  MUX21X1 U5114 ( .IN1(n6003), .IN2(n5723), .S(n5733), .Q(n6004) );
  MUX41X1 U5115 ( .IN1(n6004), .IN3(n6001), .IN2(n6002), .IN4(n4426), .S0(
        n5795), .S1(n5748), .Q(n6005) );
  MUX21X1 U5116 ( .IN1(N1764), .IN2(n509), .S(n5771), .Q(n6006) );
  MUX21X1 U5117 ( .IN1(N4510), .IN2(N4543), .S(n5771), .Q(n6007) );
  MUX21X1 U5118 ( .IN1(N1797), .IN2(N1829), .S(n5771), .Q(n6008) );
  MUX41X1 U5119 ( .IN1(n5995), .IN3(n6006), .IN2(n6008), .IN4(n6007), .S0(
        n5750), .S1(n5730), .Q(n6009) );
  MUX21X1 U5120 ( .IN1(n6010), .IN2(n6009), .S(n5788), .Q(n6012) );
  MUX41X1 U5121 ( .IN1(N1829), .IN3(N1764), .IN2(N4740), .IN4(N4773), .S0(
        n5744), .S1(n5754), .Q(n6013) );
  MUX21X1 U5122 ( .IN1(n6007), .IN2(N4549), .S(n5733), .Q(n6014) );
  MUX21X1 U5123 ( .IN1(N4909), .IN2(N4977), .S(n5771), .Q(n6015) );
  AND2X1 U5124 ( .IN1(N5010), .IN2(n5778), .Q(n6016) );
  MUX21X1 U5125 ( .IN1(n6015), .IN2(n6016), .S(n5733), .Q(n6017) );
  MUX21X1 U5126 ( .IN1(n509), .IN2(N1764), .S(n5733), .Q(n6018) );
  MUX21X1 U5127 ( .IN1(n396), .IN2(n6018), .S(n5771), .Q(n6019) );
  MUX41X1 U5128 ( .IN1(n6019), .IN3(n6014), .IN2(n6017), .IN4(n6013), .S0(
        n5795), .S1(n5747), .Q(n6020) );
  MUX41X1 U5129 ( .IN1(n6020), .IN3(n6012), .IN2(n6005), .IN4(n5999), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5651) );
  MUX21X1 U5130 ( .IN1(N4807), .IN2(N4876), .S(n5771), .Q(n6021) );
  MUX21X1 U5131 ( .IN1(N1765), .IN2(n6021), .S(n5736), .Q(n6022) );
  MUX21X1 U5132 ( .IN1(N4609), .IN2(N1765), .S(n5771), .Q(n6023) );
  MUX21X1 U5133 ( .IN1(n508), .IN2(N1765), .S(n5771), .Q(n6024) );
  MUX21X1 U5134 ( .IN1(N4352), .IN2(ID_imm_offset[10]), .S(n5771), .Q(n6025)
         );
  MUX41X1 U5135 ( .IN1(n6025), .IN3(N5290), .IN2(n6024), .IN4(n6023), .S0(
        n5750), .S1(n5729), .Q(n6026) );
  MUX21X1 U5136 ( .IN1(n6026), .IN2(n6022), .S(n5789), .Q(n6027) );
  MUX21X1 U5137 ( .IN1(N4741), .IN2(N4774), .S(n5733), .Q(n6028) );
  MUX21X1 U5138 ( .IN1(n6028), .IN2(N1765), .S(n5771), .Q(n6029) );
  MUX21X1 U5139 ( .IN1(n508), .IN2(N5225), .S(n5733), .Q(n6030) );
  MUX21X1 U5140 ( .IN1(N3015), .IN2(N4140), .S(n5771), .Q(n6031) );
  MUX21X1 U5141 ( .IN1(n6031), .IN2(n5723), .S(n5733), .Q(n6032) );
  MUX41X1 U5142 ( .IN1(n6032), .IN3(n6029), .IN2(n6030), .IN4(n4425), .S0(
        n5795), .S1(n5748), .Q(n6033) );
  MUX21X1 U5143 ( .IN1(N1765), .IN2(n508), .S(n5772), .Q(n6034) );
  MUX21X1 U5144 ( .IN1(N4511), .IN2(N4544), .S(n5772), .Q(n6035) );
  MUX21X1 U5145 ( .IN1(N1798), .IN2(N1830), .S(n5772), .Q(n6036) );
  MUX41X1 U5146 ( .IN1(n6023), .IN3(n6034), .IN2(n6036), .IN4(n6035), .S0(
        n5750), .S1(n5727), .Q(n6037) );
  MUX21X1 U5147 ( .IN1(n6038), .IN2(n6037), .S(n5789), .Q(n6040) );
  MUX41X1 U5148 ( .IN1(N1830), .IN3(N1765), .IN2(N4741), .IN4(N4774), .S0(
        n5695), .S1(n5756), .Q(n6041) );
  MUX21X1 U5149 ( .IN1(n6035), .IN2(N4548), .S(n5733), .Q(n6042) );
  MUX21X1 U5150 ( .IN1(N4910), .IN2(N4978), .S(n5772), .Q(n6043) );
  AND2X1 U5151 ( .IN1(N5011), .IN2(n5779), .Q(n6044) );
  MUX21X1 U5152 ( .IN1(n6043), .IN2(n6044), .S(n5733), .Q(n6045) );
  MUX21X1 U5153 ( .IN1(n508), .IN2(N1765), .S(n5733), .Q(n6046) );
  MUX21X1 U5154 ( .IN1(n395), .IN2(n6046), .S(n5772), .Q(n6047) );
  MUX41X1 U5155 ( .IN1(n6047), .IN3(n6042), .IN2(n6045), .IN4(n6041), .S0(
        n5795), .S1(n5748), .Q(n6048) );
  MUX41X1 U5156 ( .IN1(n6048), .IN3(n6040), .IN2(n6033), .IN4(n6027), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5652) );
  MUX21X1 U5157 ( .IN1(N4808), .IN2(N4877), .S(n5772), .Q(n6049) );
  MUX21X1 U5158 ( .IN1(N1766), .IN2(n6049), .S(n5733), .Q(n6050) );
  MUX21X1 U5159 ( .IN1(N4610), .IN2(N1766), .S(n5776), .Q(n6051) );
  MUX21X1 U5160 ( .IN1(n507), .IN2(N1766), .S(n5775), .Q(n6052) );
  MUX21X1 U5161 ( .IN1(N4351), .IN2(ID_imm_offset[10]), .S(n5775), .Q(n6053)
         );
  MUX41X1 U5162 ( .IN1(n6053), .IN3(N5291), .IN2(n6052), .IN4(n6051), .S0(
        n5750), .S1(n5726), .Q(n6054) );
  MUX21X1 U5163 ( .IN1(n6054), .IN2(n6050), .S(n5789), .Q(n6055) );
  MUX21X1 U5164 ( .IN1(N4742), .IN2(N4775), .S(n5732), .Q(n6056) );
  MUX21X1 U5165 ( .IN1(n6056), .IN2(N1766), .S(n5775), .Q(n6057) );
  MUX21X1 U5166 ( .IN1(n507), .IN2(N5226), .S(n5732), .Q(n6058) );
  MUX21X1 U5167 ( .IN1(N3016), .IN2(N4141), .S(n5775), .Q(n6059) );
  MUX21X1 U5168 ( .IN1(n6059), .IN2(n5723), .S(n5732), .Q(n6060) );
  MUX41X1 U5169 ( .IN1(n6060), .IN3(n6057), .IN2(n6058), .IN4(n4424), .S0(
        n5795), .S1(n5748), .Q(n6061) );
  MUX21X1 U5170 ( .IN1(N1766), .IN2(n507), .S(n5775), .Q(n6062) );
  MUX21X1 U5171 ( .IN1(N4512), .IN2(N4545), .S(n5775), .Q(n6063) );
  MUX21X1 U5172 ( .IN1(N1799), .IN2(N1831), .S(n5775), .Q(n6064) );
  MUX41X1 U5173 ( .IN1(n6051), .IN3(n6062), .IN2(n6064), .IN4(n6063), .S0(
        n5750), .S1(n5725), .Q(n6065) );
  MUX21X1 U5174 ( .IN1(n6066), .IN2(n6065), .S(n5789), .Q(n6068) );
  MUX41X1 U5175 ( .IN1(N1831), .IN3(N1766), .IN2(N4742), .IN4(N4775), .S0(
        n5744), .S1(n5754), .Q(n6069) );
  MUX21X1 U5176 ( .IN1(n6063), .IN2(N4547), .S(n5732), .Q(n6070) );
  MUX21X1 U5177 ( .IN1(N4911), .IN2(N4979), .S(n5775), .Q(n6071) );
  AND2X1 U5178 ( .IN1(N5012), .IN2(n5778), .Q(n6072) );
  MUX21X1 U5179 ( .IN1(n6071), .IN2(n6072), .S(n5732), .Q(n6073) );
  MUX21X1 U5180 ( .IN1(n507), .IN2(N1766), .S(n5732), .Q(n6074) );
  MUX21X1 U5181 ( .IN1(n394), .IN2(n6074), .S(n5775), .Q(n6075) );
  MUX41X1 U5182 ( .IN1(n6075), .IN3(n6070), .IN2(n6073), .IN4(n6069), .S0(
        n5795), .S1(n5749), .Q(n6076) );
  MUX41X1 U5183 ( .IN1(n6076), .IN3(n6061), .IN2(n6068), .IN4(n6055), .S0(
        ID_opcode[3]), .S1(ID_opcode[2]), .Q(N5653) );
  MUX21X1 U5184 ( .IN1(N4796), .IN2(N4865), .S(n5775), .Q(n6077) );
  MUX21X1 U5185 ( .IN1(N1754), .IN2(n6077), .S(n5732), .Q(n6078) );
  MUX21X1 U5186 ( .IN1(N4598), .IN2(N1754), .S(n5775), .Q(n6079) );
  MUX21X1 U5187 ( .IN1(n519), .IN2(N1754), .S(n5775), .Q(n6080) );
  MUX21X1 U5188 ( .IN1(N4363), .IN2(ID_imm_offset[7]), .S(n5775), .Q(n6081) );
  MUX41X1 U5189 ( .IN1(n6081), .IN3(N5279), .IN2(n6080), .IN4(n6079), .S0(
        n5751), .S1(n5724), .Q(n6082) );
  MUX21X1 U5190 ( .IN1(n6082), .IN2(n6078), .S(n5789), .Q(n6083) );
  MUX21X1 U5191 ( .IN1(N4730), .IN2(N4763), .S(n5730), .Q(n6084) );
  MUX21X1 U5192 ( .IN1(n6084), .IN2(N1754), .S(n5775), .Q(n6085) );
  MUX21X1 U5193 ( .IN1(n519), .IN2(N5214), .S(n5730), .Q(n6086) );
  MUX21X1 U5194 ( .IN1(N3004), .IN2(N4129), .S(n5775), .Q(n6087) );
  MUX21X1 U5195 ( .IN1(n6087), .IN2(n5723), .S(n5730), .Q(n6088) );
  MUX41X1 U5196 ( .IN1(n6088), .IN3(n6085), .IN2(n6086), .IN4(n4436), .S0(
        n5795), .S1(n5749), .Q(n6089) );
  MUX21X1 U5197 ( .IN1(N1754), .IN2(n519), .S(n5775), .Q(n6090) );
  MUX21X1 U5198 ( .IN1(N4500), .IN2(N4533), .S(n5775), .Q(n6091) );
  MUX21X1 U5199 ( .IN1(N1787), .IN2(N1819), .S(n5776), .Q(n6092) );
  MUX41X1 U5200 ( .IN1(n6079), .IN3(n6090), .IN2(n6092), .IN4(n6091), .S0(
        n5751), .S1(n5724), .Q(n6093) );
  MUX21X1 U5201 ( .IN1(n6094), .IN2(n6093), .S(n5789), .Q(n6096) );
  MUX41X1 U5202 ( .IN1(N1819), .IN3(N1754), .IN2(N4730), .IN4(N4763), .S0(
        n5744), .S1(n5755), .Q(n6097) );
  MUX21X1 U5203 ( .IN1(n6091), .IN2(N4559), .S(n5730), .Q(n6098) );
  MUX21X1 U5204 ( .IN1(N4899), .IN2(N4967), .S(n5776), .Q(n6099) );
  AND2X1 U5205 ( .IN1(N5000), .IN2(n5778), .Q(n6100) );
  MUX21X1 U5206 ( .IN1(n6099), .IN2(n6100), .S(n5730), .Q(n6101) );
  MUX21X1 U5207 ( .IN1(n519), .IN2(N1754), .S(n5730), .Q(n6102) );
  MUX21X1 U5208 ( .IN1(n406), .IN2(n6102), .S(n5776), .Q(n6103) );
  MUX41X1 U5209 ( .IN1(n6103), .IN3(n6098), .IN2(n6101), .IN4(n6097), .S0(
        n5795), .S1(n5749), .Q(n6104) );
  MUX41X1 U5210 ( .IN1(n6104), .IN3(n6096), .IN2(n6089), .IN4(n6083), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5641) );
  MUX21X1 U5211 ( .IN1(N4789), .IN2(N4858), .S(n5776), .Q(n6105) );
  MUX21X1 U5212 ( .IN1(N1747), .IN2(n6105), .S(n5730), .Q(n6106) );
  MUX21X1 U5213 ( .IN1(N4591), .IN2(N1747), .S(n5776), .Q(n6107) );
  MUX21X1 U5214 ( .IN1(n526), .IN2(N1747), .S(n5776), .Q(n6108) );
  MUX21X1 U5215 ( .IN1(N4370), .IN2(ID_imm_offset[0]), .S(n5776), .Q(n6109) );
  MUX41X1 U5216 ( .IN1(n6109), .IN3(N5272), .IN2(n6108), .IN4(n6107), .S0(
        n5751), .S1(n5727), .Q(n6110) );
  MUX21X1 U5217 ( .IN1(n6110), .IN2(n6106), .S(n5790), .Q(n6111) );
  MUX21X1 U5218 ( .IN1(N4723), .IN2(N4756), .S(n5730), .Q(n6112) );
  MUX21X1 U5219 ( .IN1(n6112), .IN2(N1747), .S(n5776), .Q(n6113) );
  MUX21X1 U5220 ( .IN1(n526), .IN2(N5207), .S(n5730), .Q(n6114) );
  MUX21X1 U5221 ( .IN1(N2997), .IN2(N4122), .S(n5776), .Q(n6115) );
  MUX21X1 U5222 ( .IN1(n6115), .IN2(n5723), .S(n5730), .Q(n6116) );
  MUX41X1 U5223 ( .IN1(n6116), .IN3(n6113), .IN2(n6114), .IN4(n4443), .S0(
        n5795), .S1(n5748), .Q(n6117) );
  MUX21X1 U5224 ( .IN1(N1747), .IN2(n526), .S(n5776), .Q(n6118) );
  MUX21X1 U5225 ( .IN1(N4493), .IN2(N4526), .S(n5776), .Q(n6119) );
  MUX21X1 U5226 ( .IN1(N1780), .IN2(N1812), .S(n5776), .Q(n6120) );
  MUX41X1 U5227 ( .IN1(n6107), .IN3(n6118), .IN2(n6120), .IN4(n6119), .S0(
        n5751), .S1(n5729), .Q(n6121) );
  MUX21X1 U5228 ( .IN1(n6122), .IN2(n6121), .S(n5790), .Q(n6124) );
  MUX41X1 U5229 ( .IN1(N1812), .IN3(N1747), .IN2(N4723), .IN4(N4756), .S0(
        n5744), .S1(n5756), .Q(n6125) );
  MUX21X1 U5230 ( .IN1(n6119), .IN2(N4566), .S(n5730), .Q(n6126) );
  MUX21X1 U5231 ( .IN1(N4892), .IN2(N4960), .S(n5776), .Q(n6127) );
  AND2X1 U5232 ( .IN1(N4993), .IN2(n5779), .Q(n6128) );
  MUX21X1 U5233 ( .IN1(n6127), .IN2(n6128), .S(n5730), .Q(n6129) );
  MUX21X1 U5234 ( .IN1(n526), .IN2(N1747), .S(n5730), .Q(n6130) );
  MUX21X1 U5235 ( .IN1(n413), .IN2(n6130), .S(n5776), .Q(n6131) );
  MUX41X1 U5236 ( .IN1(n6131), .IN3(n6126), .IN2(n6129), .IN4(n6125), .S0(
        n5795), .S1(n5749), .Q(n6132) );
  MUX41X1 U5237 ( .IN1(n6132), .IN3(n6124), .IN2(n6117), .IN4(n6111), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5634) );
  MUX21X1 U5238 ( .IN1(N4790), .IN2(N4859), .S(n5776), .Q(n6133) );
  MUX21X1 U5239 ( .IN1(N1748), .IN2(n6133), .S(n5731), .Q(n6134) );
  MUX21X1 U5240 ( .IN1(N4592), .IN2(N1748), .S(n5774), .Q(n6135) );
  MUX21X1 U5241 ( .IN1(n525), .IN2(N1748), .S(n5774), .Q(n6136) );
  MUX21X1 U5242 ( .IN1(N4369), .IN2(ID_imm_offset[1]), .S(n5774), .Q(n6137) );
  MUX41X1 U5243 ( .IN1(n6137), .IN3(N5273), .IN2(n6136), .IN4(n6135), .S0(
        n5751), .S1(n5729), .Q(n6138) );
  MUX21X1 U5244 ( .IN1(n6138), .IN2(n6134), .S(n5789), .Q(n6139) );
  MUX21X1 U5245 ( .IN1(N4724), .IN2(N4757), .S(n5731), .Q(n6140) );
  MUX21X1 U5246 ( .IN1(n6140), .IN2(N1748), .S(n5774), .Q(n6141) );
  MUX21X1 U5247 ( .IN1(n525), .IN2(N5208), .S(n5731), .Q(n6142) );
  MUX21X1 U5248 ( .IN1(N2998), .IN2(N4123), .S(n5774), .Q(n6143) );
  MUX21X1 U5249 ( .IN1(n6143), .IN2(n5723), .S(n5731), .Q(n6144) );
  MUX41X1 U5250 ( .IN1(n6144), .IN3(n6141), .IN2(n6142), .IN4(n4442), .S0(
        n5795), .S1(n5749), .Q(n6145) );
  MUX21X1 U5251 ( .IN1(N1748), .IN2(n525), .S(n5774), .Q(n6146) );
  MUX21X1 U5252 ( .IN1(N4494), .IN2(N4527), .S(n5774), .Q(n6147) );
  MUX21X1 U5253 ( .IN1(N1781), .IN2(N1813), .S(n5774), .Q(n6148) );
  MUX41X1 U5254 ( .IN1(n6135), .IN3(n6146), .IN2(n6148), .IN4(n6147), .S0(
        n5751), .S1(n5729), .Q(n6149) );
  MUX21X1 U5255 ( .IN1(n6150), .IN2(n6149), .S(n5789), .Q(n6152) );
  MUX41X1 U5256 ( .IN1(N1813), .IN3(N1748), .IN2(N4724), .IN4(N4757), .S0(
        n5743), .S1(n5755), .Q(n6153) );
  MUX21X1 U5257 ( .IN1(n6147), .IN2(N4565), .S(n5731), .Q(n6154) );
  MUX21X1 U5258 ( .IN1(N4893), .IN2(N4961), .S(n5774), .Q(n6155) );
  AND2X1 U5259 ( .IN1(N4994), .IN2(n5778), .Q(n6156) );
  MUX21X1 U5260 ( .IN1(n6155), .IN2(n6156), .S(n5731), .Q(n6157) );
  MUX21X1 U5261 ( .IN1(n525), .IN2(N1748), .S(n5731), .Q(n6158) );
  MUX21X1 U5262 ( .IN1(n412), .IN2(n6158), .S(n5774), .Q(n6159) );
  MUX41X1 U5263 ( .IN1(n6159), .IN3(n6154), .IN2(n6157), .IN4(n6153), .S0(
        n5794), .S1(n5749), .Q(n6160) );
  MUX41X1 U5264 ( .IN1(n6160), .IN3(n6152), .IN2(n6145), .IN4(n6139), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5635) );
  MUX21X1 U5265 ( .IN1(N4791), .IN2(N4860), .S(n5774), .Q(n6161) );
  MUX21X1 U5266 ( .IN1(N1749), .IN2(n6161), .S(n5731), .Q(n6162) );
  MUX21X1 U5267 ( .IN1(N4593), .IN2(N1749), .S(n5774), .Q(n6163) );
  MUX21X1 U5268 ( .IN1(n524), .IN2(N1749), .S(n5774), .Q(n6164) );
  MUX21X1 U5269 ( .IN1(N4368), .IN2(ID_imm_offset[2]), .S(n5774), .Q(n6165) );
  MUX41X1 U5270 ( .IN1(n6165), .IN3(N5274), .IN2(n6164), .IN4(n6163), .S0(
        n5751), .S1(n5728), .Q(n6166) );
  MUX21X1 U5271 ( .IN1(n6166), .IN2(n6162), .S(n5790), .Q(n6167) );
  MUX21X1 U5272 ( .IN1(N4725), .IN2(N4758), .S(n5731), .Q(n6168) );
  MUX21X1 U5273 ( .IN1(n6168), .IN2(N1749), .S(n5774), .Q(n6169) );
  MUX21X1 U5274 ( .IN1(n524), .IN2(N5209), .S(n5731), .Q(n6170) );
  MUX21X1 U5275 ( .IN1(N2999), .IN2(N4124), .S(n5774), .Q(n6171) );
  MUX21X1 U5276 ( .IN1(n6171), .IN2(n5723), .S(n5731), .Q(n6172) );
  MUX41X1 U5277 ( .IN1(n6172), .IN3(n6169), .IN2(n6170), .IN4(n4441), .S0(
        n5794), .S1(n5749), .Q(n6173) );
  MUX21X1 U5278 ( .IN1(N1749), .IN2(n524), .S(n5774), .Q(n6174) );
  MUX21X1 U5279 ( .IN1(N4495), .IN2(N4528), .S(n5774), .Q(n6175) );
  MUX21X1 U5280 ( .IN1(N1782), .IN2(N1814), .S(n5773), .Q(n6176) );
  MUX41X1 U5281 ( .IN1(n6163), .IN3(n6174), .IN2(n6176), .IN4(n6175), .S0(
        n5751), .S1(n5726), .Q(n6177) );
  MUX21X1 U5282 ( .IN1(n6178), .IN2(n6177), .S(n5790), .Q(n6180) );
  MUX41X1 U5283 ( .IN1(N1814), .IN3(N1749), .IN2(N4725), .IN4(N4758), .S0(
        n5744), .S1(n5755), .Q(n6181) );
  MUX21X1 U5284 ( .IN1(n6175), .IN2(N4564), .S(n5731), .Q(n6182) );
  MUX21X1 U5285 ( .IN1(N4894), .IN2(N4962), .S(n5773), .Q(n6183) );
  AND2X1 U5286 ( .IN1(N4995), .IN2(n5778), .Q(n6184) );
  MUX21X1 U5287 ( .IN1(n6183), .IN2(n6184), .S(n5731), .Q(n6185) );
  MUX21X1 U5288 ( .IN1(n524), .IN2(N1749), .S(n5731), .Q(n6186) );
  MUX21X1 U5289 ( .IN1(n411), .IN2(n6186), .S(n5773), .Q(n6187) );
  MUX41X1 U5290 ( .IN1(n6187), .IN3(n6182), .IN2(n6185), .IN4(n6181), .S0(
        n5794), .S1(n5748), .Q(n6188) );
  MUX41X1 U5291 ( .IN1(n6188), .IN3(n6180), .IN2(n6173), .IN4(n6167), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5636) );
  MUX21X1 U5292 ( .IN1(N4792), .IN2(N4861), .S(n5773), .Q(n6189) );
  MUX21X1 U5293 ( .IN1(N1750), .IN2(n6189), .S(n5731), .Q(n6190) );
  MUX21X1 U5294 ( .IN1(N4594), .IN2(N1750), .S(n5773), .Q(n6191) );
  MUX21X1 U5295 ( .IN1(n523), .IN2(N1750), .S(n5773), .Q(n6192) );
  MUX21X1 U5296 ( .IN1(N4367), .IN2(ID_imm_offset[3]), .S(n5773), .Q(n6193) );
  MUX41X1 U5297 ( .IN1(n6193), .IN3(N5275), .IN2(n6192), .IN4(n6191), .S0(
        n5751), .S1(n5725), .Q(n6194) );
  MUX21X1 U5298 ( .IN1(n6194), .IN2(n6190), .S(n5789), .Q(n6195) );
  MUX21X1 U5299 ( .IN1(N4726), .IN2(N4759), .S(n5731), .Q(n6196) );
  MUX21X1 U5300 ( .IN1(n6196), .IN2(N1750), .S(n5773), .Q(n6197) );
  MUX21X1 U5301 ( .IN1(n523), .IN2(N5210), .S(n5731), .Q(n6198) );
  MUX21X1 U5302 ( .IN1(N3000), .IN2(N4125), .S(n5773), .Q(n6199) );
  MUX21X1 U5303 ( .IN1(n6199), .IN2(n5723), .S(n5731), .Q(n6200) );
  MUX41X1 U5304 ( .IN1(n6200), .IN3(n6197), .IN2(n6198), .IN4(n4440), .S0(
        n5794), .S1(n5750), .Q(n6201) );
  MUX21X1 U5305 ( .IN1(N1750), .IN2(n523), .S(n5773), .Q(n6202) );
  MUX21X1 U5306 ( .IN1(N4496), .IN2(N4529), .S(n5773), .Q(n6203) );
  MUX21X1 U5307 ( .IN1(N1783), .IN2(N1815), .S(n5773), .Q(n6204) );
  MUX41X1 U5308 ( .IN1(n6191), .IN3(n6202), .IN2(n6204), .IN4(n6203), .S0(
        n5751), .S1(n5725), .Q(n6205) );
  MUX21X1 U5309 ( .IN1(n6206), .IN2(n6205), .S(n5791), .Q(n6208) );
  MUX41X1 U5310 ( .IN1(N1815), .IN3(N1750), .IN2(N4726), .IN4(N4759), .S0(
        n5744), .S1(n5755), .Q(n6209) );
  MUX21X1 U5311 ( .IN1(n6203), .IN2(N4563), .S(n5732), .Q(n6210) );
  MUX21X1 U5312 ( .IN1(N4895), .IN2(N4963), .S(n5773), .Q(n6211) );
  AND2X1 U5313 ( .IN1(N4996), .IN2(n5778), .Q(n6212) );
  MUX21X1 U5314 ( .IN1(n6211), .IN2(n6212), .S(n5732), .Q(n6213) );
  MUX21X1 U5315 ( .IN1(n523), .IN2(N1750), .S(n5732), .Q(n6214) );
  MUX21X1 U5316 ( .IN1(n410), .IN2(n6214), .S(n5773), .Q(n6215) );
  MUX41X1 U5317 ( .IN1(n6215), .IN3(n6210), .IN2(n6213), .IN4(n6209), .S0(
        n5794), .S1(n5750), .Q(n6216) );
  MUX41X1 U5318 ( .IN1(n6216), .IN3(n6208), .IN2(n6201), .IN4(n6195), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5637) );
  MUX21X1 U5319 ( .IN1(N4793), .IN2(N4862), .S(n5775), .Q(n6217) );
  MUX21X1 U5320 ( .IN1(N1751), .IN2(n6217), .S(n5732), .Q(n6218) );
  MUX21X1 U5321 ( .IN1(N4595), .IN2(N1751), .S(n5773), .Q(n6219) );
  MUX21X1 U5322 ( .IN1(n522), .IN2(N1751), .S(n5773), .Q(n6220) );
  MUX21X1 U5323 ( .IN1(N4366), .IN2(ID_imm_offset[4]), .S(n5773), .Q(n6221) );
  MUX41X1 U5324 ( .IN1(n6221), .IN3(N5276), .IN2(n6220), .IN4(n6219), .S0(
        n5751), .S1(n5725), .Q(n6222) );
  MUX21X1 U5325 ( .IN1(n6222), .IN2(n6218), .S(n5790), .Q(n6223) );
  MUX21X1 U5326 ( .IN1(N4727), .IN2(N4760), .S(n5732), .Q(n6224) );
  MUX21X1 U5327 ( .IN1(n6224), .IN2(N1751), .S(n5772), .Q(n6225) );
  MUX21X1 U5328 ( .IN1(n522), .IN2(N5211), .S(n5732), .Q(n6226) );
  MUX21X1 U5329 ( .IN1(N3001), .IN2(N4126), .S(n5772), .Q(n6227) );
  MUX21X1 U5330 ( .IN1(n6227), .IN2(n5723), .S(n5732), .Q(n6228) );
  MUX41X1 U5331 ( .IN1(n6228), .IN3(n6225), .IN2(n6226), .IN4(n4439), .S0(
        n5794), .S1(n5750), .Q(n6229) );
  MUX21X1 U5332 ( .IN1(N1751), .IN2(n522), .S(n5772), .Q(n6230) );
  MUX21X1 U5333 ( .IN1(N4497), .IN2(N4530), .S(n5772), .Q(n6231) );
  MUX21X1 U5334 ( .IN1(N1784), .IN2(N1816), .S(n5772), .Q(n6232) );
  MUX41X1 U5335 ( .IN1(n6219), .IN3(n6230), .IN2(n6232), .IN4(n6231), .S0(
        n5751), .S1(n5724), .Q(n6233) );
  MUX21X1 U5336 ( .IN1(n6234), .IN2(n6233), .S(n5791), .Q(n6236) );
  MUX41X1 U5337 ( .IN1(N1816), .IN3(N1751), .IN2(N4727), .IN4(N4760), .S0(
        n5695), .S1(n5754), .Q(n6237) );
  MUX21X1 U5338 ( .IN1(n6231), .IN2(N4562), .S(n5732), .Q(n6238) );
  MUX21X1 U5339 ( .IN1(N4896), .IN2(N4964), .S(n5772), .Q(n6239) );
  AND2X1 U5340 ( .IN1(N4997), .IN2(n5779), .Q(n6240) );
  MUX21X1 U5341 ( .IN1(n6239), .IN2(n6240), .S(n5732), .Q(n6241) );
  MUX21X1 U5342 ( .IN1(n522), .IN2(N1751), .S(n5732), .Q(n6242) );
  MUX21X1 U5343 ( .IN1(n409), .IN2(n6242), .S(n5772), .Q(n6243) );
  MUX41X1 U5344 ( .IN1(n6243), .IN3(n6238), .IN2(n6241), .IN4(n6237), .S0(
        n5794), .S1(n5750), .Q(n6244) );
  MUX41X1 U5345 ( .IN1(n6244), .IN3(n6236), .IN2(n6229), .IN4(n6223), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5638) );
  MUX21X1 U5346 ( .IN1(N4794), .IN2(N4863), .S(n5772), .Q(n6245) );
  MUX21X1 U5347 ( .IN1(N1752), .IN2(n6245), .S(n5730), .Q(n6246) );
  MUX21X1 U5348 ( .IN1(N4596), .IN2(N1752), .S(n5772), .Q(n6247) );
  MUX21X1 U5349 ( .IN1(n521), .IN2(N1752), .S(n5772), .Q(n6248) );
  MUX21X1 U5350 ( .IN1(N4365), .IN2(ID_imm_offset[5]), .S(n5772), .Q(n6249) );
  MUX41X1 U5351 ( .IN1(n6249), .IN3(N5277), .IN2(n6248), .IN4(n6247), .S0(
        n5751), .S1(n5724), .Q(n6250) );
  MUX21X1 U5352 ( .IN1(n6250), .IN2(n6246), .S(n5791), .Q(n6251) );
  MUX21X1 U5353 ( .IN1(N4728), .IN2(N4761), .S(n5732), .Q(n6252) );
  MUX21X1 U5354 ( .IN1(n6252), .IN2(N1752), .S(n5773), .Q(n6253) );
  MUX21X1 U5355 ( .IN1(n521), .IN2(N5212), .S(n5742), .Q(n6254) );
  MUX21X1 U5356 ( .IN1(N3002), .IN2(N4127), .S(n5761), .Q(n6255) );
  MUX21X1 U5357 ( .IN1(n6255), .IN2(n5723), .S(n5740), .Q(n6256) );
  MUX41X1 U5358 ( .IN1(n6256), .IN3(n6253), .IN2(n6254), .IN4(n4438), .S0(
        n5794), .S1(n5749), .Q(n6257) );
  MUX21X1 U5359 ( .IN1(N1752), .IN2(n521), .S(n5761), .Q(n6258) );
  MUX21X1 U5360 ( .IN1(N4498), .IN2(N4531), .S(n5761), .Q(n6259) );
  MUX21X1 U5361 ( .IN1(N1785), .IN2(N1817), .S(n5761), .Q(n6260) );
  MUX41X1 U5362 ( .IN1(n6247), .IN3(n6258), .IN2(n6260), .IN4(n6259), .S0(
        n5751), .S1(n5724), .Q(n6261) );
  MUX21X1 U5363 ( .IN1(n6262), .IN2(n6261), .S(n5790), .Q(n6264) );
  MUX41X1 U5364 ( .IN1(N1817), .IN3(N1752), .IN2(N4728), .IN4(N4761), .S0(
        n5695), .S1(n5754), .Q(n6265) );
  MUX21X1 U5365 ( .IN1(n6259), .IN2(N4561), .S(n5740), .Q(n6266) );
  MUX21X1 U5366 ( .IN1(N4897), .IN2(N4965), .S(n5761), .Q(n6267) );
  AND2X1 U5367 ( .IN1(N4998), .IN2(n5779), .Q(n6268) );
  MUX21X1 U5368 ( .IN1(n6267), .IN2(n6268), .S(n5740), .Q(n6269) );
  MUX21X1 U5369 ( .IN1(n521), .IN2(N1752), .S(n5740), .Q(n6270) );
  MUX21X1 U5370 ( .IN1(n408), .IN2(n6270), .S(n5761), .Q(n6271) );
  MUX41X1 U5371 ( .IN1(n6271), .IN3(n6266), .IN2(n6269), .IN4(n6265), .S0(
        n5794), .S1(n5748), .Q(n6272) );
  MUX41X1 U5372 ( .IN1(n6272), .IN3(n6264), .IN2(n6257), .IN4(n6251), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5639) );
  MUX21X1 U5373 ( .IN1(N4795), .IN2(N4864), .S(n5761), .Q(n6273) );
  MUX21X1 U5374 ( .IN1(N1753), .IN2(n6273), .S(n5740), .Q(n6274) );
  MUX21X1 U5375 ( .IN1(N4597), .IN2(N1753), .S(n5761), .Q(n6275) );
  MUX21X1 U5376 ( .IN1(n520), .IN2(N1753), .S(n5760), .Q(n6276) );
  MUX21X1 U5377 ( .IN1(N4364), .IN2(ID_imm_offset[6]), .S(n5760), .Q(n6277) );
  MUX41X1 U5378 ( .IN1(n6277), .IN3(N5278), .IN2(n6276), .IN4(n6275), .S0(
        n5752), .S1(n5724), .Q(n6278) );
  MUX21X1 U5379 ( .IN1(n6278), .IN2(n6274), .S(n5791), .Q(n6279) );
  MUX21X1 U5380 ( .IN1(N4729), .IN2(N4762), .S(n5740), .Q(n6280) );
  MUX21X1 U5381 ( .IN1(n6280), .IN2(N1753), .S(n5760), .Q(n6281) );
  MUX21X1 U5382 ( .IN1(n520), .IN2(N5213), .S(n5740), .Q(n6282) );
  MUX21X1 U5383 ( .IN1(N3003), .IN2(N4128), .S(n5760), .Q(n6283) );
  MUX21X1 U5384 ( .IN1(n6283), .IN2(n5723), .S(n5741), .Q(n6284) );
  MUX41X1 U5385 ( .IN1(n6284), .IN3(n6281), .IN2(n6282), .IN4(n4437), .S0(
        n5794), .S1(n5749), .Q(n6285) );
  MUX21X1 U5386 ( .IN1(N1753), .IN2(n520), .S(n5760), .Q(n6286) );
  MUX21X1 U5387 ( .IN1(N4499), .IN2(N4532), .S(n5760), .Q(n6287) );
  MUX21X1 U5388 ( .IN1(N1786), .IN2(N1818), .S(n5760), .Q(n6288) );
  MUX41X1 U5389 ( .IN1(n6275), .IN3(n6286), .IN2(n6288), .IN4(n6287), .S0(
        n5751), .S1(n5724), .Q(n6289) );
  MUX21X1 U5390 ( .IN1(n6290), .IN2(n6289), .S(n5790), .Q(n6292) );
  MUX41X1 U5391 ( .IN1(N1818), .IN3(N1753), .IN2(N4729), .IN4(N4762), .S0(
        n5744), .S1(n5754), .Q(n6293) );
  MUX21X1 U5392 ( .IN1(n6287), .IN2(N4560), .S(n5741), .Q(n6294) );
  MUX21X1 U5393 ( .IN1(N4898), .IN2(N4966), .S(n5760), .Q(n6295) );
  AND2X1 U5394 ( .IN1(N4999), .IN2(n5779), .Q(n6296) );
  MUX21X1 U5395 ( .IN1(n6295), .IN2(n6296), .S(n5741), .Q(n6297) );
  MUX21X1 U5396 ( .IN1(n520), .IN2(N1753), .S(n5741), .Q(n6298) );
  MUX21X1 U5397 ( .IN1(n407), .IN2(n6298), .S(n5760), .Q(n6299) );
  MUX41X1 U5398 ( .IN1(n6299), .IN3(n6294), .IN2(n6297), .IN4(n6293), .S0(
        n5794), .S1(n5749), .Q(n6300) );
  MUX41X1 U5399 ( .IN1(n6300), .IN3(n6292), .IN2(n6285), .IN4(n6279), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5640) );
  MUX21X1 U5400 ( .IN1(N4797), .IN2(N4866), .S(n5760), .Q(n6301) );
  MUX21X1 U5401 ( .IN1(N1755), .IN2(n6301), .S(n5741), .Q(n6302) );
  MUX21X1 U5402 ( .IN1(N4599), .IN2(N1755), .S(n5760), .Q(n6303) );
  MUX21X1 U5403 ( .IN1(n518), .IN2(N1755), .S(n5760), .Q(n6304) );
  MUX21X1 U5404 ( .IN1(N4362), .IN2(ID_imm_offset[8]), .S(n5760), .Q(n6305) );
  MUX41X1 U5405 ( .IN1(n6305), .IN3(N5280), .IN2(n6304), .IN4(n6303), .S0(
        n5752), .S1(n5725), .Q(n6306) );
  MUX21X1 U5406 ( .IN1(n6306), .IN2(n6302), .S(n5791), .Q(n6307) );
  MUX21X1 U5407 ( .IN1(N4731), .IN2(N4764), .S(n5741), .Q(n6308) );
  MUX21X1 U5408 ( .IN1(n6308), .IN2(N1755), .S(n5760), .Q(n6309) );
  MUX21X1 U5409 ( .IN1(n518), .IN2(N5215), .S(n5741), .Q(n6310) );
  MUX21X1 U5410 ( .IN1(N3005), .IN2(N4130), .S(n5760), .Q(n6311) );
  MUX21X1 U5411 ( .IN1(n6311), .IN2(n5723), .S(n5741), .Q(n6312) );
  MUX41X1 U5412 ( .IN1(n6312), .IN3(n6309), .IN2(n6310), .IN4(n4435), .S0(
        n5794), .S1(n5749), .Q(n6313) );
  MUX21X1 U5413 ( .IN1(N1755), .IN2(n518), .S(n5760), .Q(n6314) );
  MUX21X1 U5414 ( .IN1(N4501), .IN2(N4534), .S(n5760), .Q(n6315) );
  MUX21X1 U5415 ( .IN1(N1788), .IN2(N1820), .S(n5760), .Q(n6316) );
  MUX41X1 U5416 ( .IN1(n6303), .IN3(n6314), .IN2(n6316), .IN4(n6315), .S0(
        n5751), .S1(n5725), .Q(n6317) );
  MUX21X1 U5417 ( .IN1(n6318), .IN2(n6317), .S(n5791), .Q(n6320) );
  MUX41X1 U5418 ( .IN1(N1820), .IN3(N1755), .IN2(N4731), .IN4(N4764), .S0(
        n5744), .S1(n5755), .Q(n6321) );
  MUX21X1 U5419 ( .IN1(n6315), .IN2(N4558), .S(n5741), .Q(n6322) );
  MUX21X1 U5420 ( .IN1(N4900), .IN2(N4968), .S(n5759), .Q(n6323) );
  AND2X1 U5421 ( .IN1(N5001), .IN2(n5779), .Q(n6324) );
  MUX21X1 U5422 ( .IN1(n6323), .IN2(n6324), .S(n5741), .Q(n6325) );
  MUX21X1 U5423 ( .IN1(n518), .IN2(N1755), .S(n5741), .Q(n6326) );
  MUX21X1 U5424 ( .IN1(n405), .IN2(n6326), .S(n5759), .Q(n6327) );
  MUX41X1 U5425 ( .IN1(n6327), .IN3(n6322), .IN2(n6325), .IN4(n6321), .S0(
        n5794), .S1(n5749), .Q(n6328) );
  MUX41X1 U5426 ( .IN1(n6328), .IN3(n6320), .IN2(n6313), .IN4(n6307), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5642) );
  MUX21X1 U5427 ( .IN1(N4798), .IN2(N4867), .S(n5759), .Q(n6329) );
  MUX21X1 U5428 ( .IN1(N1756), .IN2(n6329), .S(n5741), .Q(n6330) );
  MUX21X1 U5429 ( .IN1(N4600), .IN2(N1756), .S(n5759), .Q(n6331) );
  MUX21X1 U5430 ( .IN1(n517), .IN2(N1756), .S(n5759), .Q(n6332) );
  MUX21X1 U5431 ( .IN1(N4361), .IN2(ID_imm_offset[9]), .S(n5759), .Q(n6333) );
  MUX41X1 U5432 ( .IN1(n6333), .IN3(N5281), .IN2(n6332), .IN4(n6331), .S0(
        n5752), .S1(n5727), .Q(n6334) );
  MUX21X1 U5433 ( .IN1(n6334), .IN2(n6330), .S(n5791), .Q(n6335) );
  MUX21X1 U5434 ( .IN1(N4732), .IN2(N4765), .S(n5741), .Q(n6336) );
  MUX21X1 U5435 ( .IN1(n6336), .IN2(N1756), .S(n5759), .Q(n6337) );
  MUX21X1 U5436 ( .IN1(n517), .IN2(N5216), .S(n5741), .Q(n6338) );
  MUX21X1 U5437 ( .IN1(N3006), .IN2(N4131), .S(n5759), .Q(n6339) );
  MUX21X1 U5438 ( .IN1(n6339), .IN2(n5723), .S(n5741), .Q(n6340) );
  MUX41X1 U5439 ( .IN1(n6340), .IN3(n6337), .IN2(n6338), .IN4(n4434), .S0(
        n5794), .S1(n5748), .Q(n6341) );
  MUX21X1 U5440 ( .IN1(N1756), .IN2(n517), .S(n5759), .Q(n6342) );
  MUX21X1 U5441 ( .IN1(N4502), .IN2(N4535), .S(n5759), .Q(n6343) );
  MUX21X1 U5442 ( .IN1(N1789), .IN2(N1821), .S(n5759), .Q(n6344) );
  MUX41X1 U5443 ( .IN1(n6331), .IN3(n6342), .IN2(n6344), .IN4(n6343), .S0(
        n5752), .S1(n5726), .Q(n6345) );
  MUX21X1 U5444 ( .IN1(n6346), .IN2(n6345), .S(n5791), .Q(n6348) );
  MUX41X1 U5445 ( .IN1(N1821), .IN3(N1756), .IN2(N4732), .IN4(N4765), .S0(
        n5744), .S1(n5755), .Q(n6349) );
  MUX21X1 U5446 ( .IN1(n6343), .IN2(N4557), .S(n5741), .Q(n6350) );
  MUX21X1 U5447 ( .IN1(N4901), .IN2(N4969), .S(n5759), .Q(n6351) );
  AND2X1 U5448 ( .IN1(N5002), .IN2(n5778), .Q(n6352) );
  MUX21X1 U5449 ( .IN1(n6351), .IN2(n6352), .S(n5741), .Q(n6353) );
  MUX21X1 U5450 ( .IN1(n517), .IN2(N1756), .S(n5741), .Q(n6354) );
  MUX21X1 U5451 ( .IN1(n404), .IN2(n6354), .S(n5759), .Q(n6355) );
  MUX41X1 U5452 ( .IN1(n6355), .IN3(n6350), .IN2(n6353), .IN4(n6349), .S0(
        n5794), .S1(n5748), .Q(n6356) );
  MUX41X1 U5453 ( .IN1(n6356), .IN3(n6348), .IN2(n6341), .IN4(n6335), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5643) );
  MUX21X1 U5454 ( .IN1(N4786), .IN2(N4855), .S(n5759), .Q(n6357) );
  MUX21X1 U5455 ( .IN1(N1744), .IN2(n6357), .S(n5742), .Q(n6358) );
  MUX21X1 U5456 ( .IN1(N4588), .IN2(N1744), .S(n5759), .Q(n6359) );
  MUX21X1 U5457 ( .IN1(n529), .IN2(N1744), .S(n5759), .Q(n6360) );
  AND2X1 U5458 ( .IN1(N4373), .IN2(n5786), .Q(n6361) );
  MUX41X1 U5459 ( .IN1(n6361), .IN3(N5269), .IN2(n6360), .IN4(n6359), .S0(
        n5751), .S1(n5726), .Q(n6362) );
  MUX21X1 U5460 ( .IN1(n6362), .IN2(n6358), .S(n5792), .Q(n6363) );
  MUX21X1 U5461 ( .IN1(N4720), .IN2(N4753), .S(n5742), .Q(n6364) );
  MUX21X1 U5462 ( .IN1(n6364), .IN2(N1744), .S(n5759), .Q(n6365) );
  MUX21X1 U5463 ( .IN1(n529), .IN2(N5204), .S(n5742), .Q(n6366) );
  MUX41X1 U5464 ( .IN1(N2994), .IN3(N4119), .IN2(ID_imm_offset[7]), .IN4(
        ID_imm_offset[8]), .S0(n5777), .S1(n5729), .Q(n6367) );
  MUX41X1 U5465 ( .IN1(n6367), .IN3(n6365), .IN2(n6366), .IN4(n4446), .S0(
        n5793), .S1(n5748), .Q(n6368) );
  MUX21X1 U5466 ( .IN1(N1744), .IN2(n529), .S(n5759), .Q(n6369) );
  MUX21X1 U5467 ( .IN1(N4490), .IN2(N4523), .S(n5758), .Q(n6370) );
  MUX21X1 U5468 ( .IN1(N1777), .IN2(N1809), .S(n5758), .Q(n6371) );
  MUX41X1 U5469 ( .IN1(n6359), .IN3(n6369), .IN2(n6371), .IN4(n6370), .S0(
        n5752), .S1(n5726), .Q(n6372) );
  MUX21X1 U5470 ( .IN1(n6373), .IN2(n6372), .S(n5792), .Q(n6375) );
  MUX41X1 U5471 ( .IN1(N1809), .IN3(N1744), .IN2(N4720), .IN4(N4753), .S0(
        n5743), .S1(n5756), .Q(n6376) );
  MUX21X1 U5472 ( .IN1(n6370), .IN2(N4569), .S(n5742), .Q(n6377) );
  MUX21X1 U5473 ( .IN1(N4889), .IN2(N4957), .S(n5758), .Q(n6378) );
  AND2X1 U5474 ( .IN1(N4990), .IN2(n5779), .Q(n6379) );
  MUX21X1 U5475 ( .IN1(n6378), .IN2(n6379), .S(n5742), .Q(n6380) );
  MUX21X1 U5476 ( .IN1(n529), .IN2(N1744), .S(n5742), .Q(n6381) );
  MUX21X1 U5477 ( .IN1(n416), .IN2(n6381), .S(n5758), .Q(n6382) );
  MUX41X1 U5478 ( .IN1(n6382), .IN3(n6377), .IN2(n6380), .IN4(n6376), .S0(
        n5793), .S1(n5748), .Q(n6383) );
  MUX41X1 U5479 ( .IN1(n6383), .IN3(n6375), .IN2(n6368), .IN4(n6363), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5631) );
  MUX21X1 U5480 ( .IN1(N4787), .IN2(N4856), .S(n5758), .Q(n6384) );
  MUX21X1 U5481 ( .IN1(N1745), .IN2(n6384), .S(n5742), .Q(n6385) );
  MUX21X1 U5482 ( .IN1(N4589), .IN2(N1745), .S(n5758), .Q(n6386) );
  MUX21X1 U5483 ( .IN1(n528), .IN2(N1745), .S(n5758), .Q(n6387) );
  AND2X1 U5484 ( .IN1(N4372), .IN2(n5785), .Q(n6388) );
  MUX41X1 U5485 ( .IN1(n6388), .IN3(N5270), .IN2(n6387), .IN4(n6386), .S0(
        n5752), .S1(n5728), .Q(n6389) );
  MUX21X1 U5486 ( .IN1(n6389), .IN2(n6385), .S(n5791), .Q(n6390) );
  MUX21X1 U5487 ( .IN1(N4721), .IN2(N4754), .S(n5742), .Q(n6391) );
  MUX21X1 U5488 ( .IN1(n6391), .IN2(N1745), .S(n5758), .Q(n6392) );
  MUX21X1 U5489 ( .IN1(n528), .IN2(N5205), .S(n5742), .Q(n6393) );
  MUX41X1 U5490 ( .IN1(N2995), .IN3(N4120), .IN2(ID_imm_offset[7]), .IN4(
        ID_imm_offset[9]), .S0(n5777), .S1(n5729), .Q(n6394) );
  MUX41X1 U5491 ( .IN1(n6394), .IN3(n6392), .IN2(n6393), .IN4(n4445), .S0(
        n5793), .S1(n5748), .Q(n6395) );
  MUX21X1 U5492 ( .IN1(N1745), .IN2(n528), .S(n5758), .Q(n6396) );
  MUX21X1 U5493 ( .IN1(N4491), .IN2(N4524), .S(n5758), .Q(n6397) );
  MUX21X1 U5494 ( .IN1(N1778), .IN2(N1810), .S(n5758), .Q(n6398) );
  MUX41X1 U5495 ( .IN1(n6386), .IN3(n6396), .IN2(n6398), .IN4(n6397), .S0(
        n5752), .S1(n5730), .Q(n6399) );
  MUX21X1 U5496 ( .IN1(n6400), .IN2(n6399), .S(n5792), .Q(n6402) );
  MUX41X1 U5497 ( .IN1(N1810), .IN3(N1745), .IN2(N4721), .IN4(N4754), .S0(
        n5743), .S1(n5755), .Q(n6403) );
  MUX21X1 U5498 ( .IN1(n6397), .IN2(N4568), .S(n5742), .Q(n6404) );
  MUX21X1 U5499 ( .IN1(N4890), .IN2(N4958), .S(n5758), .Q(n6405) );
  AND2X1 U5500 ( .IN1(N4991), .IN2(n5778), .Q(n6406) );
  MUX21X1 U5501 ( .IN1(n6405), .IN2(n6406), .S(n5742), .Q(n6407) );
  MUX21X1 U5502 ( .IN1(n528), .IN2(N1745), .S(n5742), .Q(n6408) );
  MUX21X1 U5503 ( .IN1(n415), .IN2(n6408), .S(n5757), .Q(n6409) );
  MUX41X1 U5504 ( .IN1(n6409), .IN3(n6404), .IN2(n6407), .IN4(n6403), .S0(
        n5793), .S1(n5747), .Q(n6410) );
  MUX41X1 U5505 ( .IN1(n6410), .IN3(n6402), .IN2(n6395), .IN4(n6390), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5632) );
  MUX21X1 U5506 ( .IN1(N4788), .IN2(N4857), .S(n5757), .Q(n6411) );
  MUX21X1 U5507 ( .IN1(N1746), .IN2(n6411), .S(n5742), .Q(n6412) );
  MUX21X1 U5508 ( .IN1(N4590), .IN2(N1746), .S(n5757), .Q(n6413) );
  MUX21X1 U5509 ( .IN1(n527), .IN2(N1746), .S(n5758), .Q(n6414) );
  AND2X1 U5510 ( .IN1(N4371), .IN2(n5786), .Q(n6415) );
  MUX41X1 U5511 ( .IN1(n6415), .IN3(N5271), .IN2(n6414), .IN4(n6413), .S0(
        n5752), .S1(n5728), .Q(n6416) );
  MUX21X1 U5512 ( .IN1(n6416), .IN2(n6412), .S(n5792), .Q(n6417) );
  MUX21X1 U5513 ( .IN1(N4722), .IN2(N4755), .S(n5743), .Q(n6418) );
  MUX21X1 U5514 ( .IN1(n6418), .IN2(N1746), .S(n5757), .Q(n6419) );
  MUX21X1 U5515 ( .IN1(n527), .IN2(N5206), .S(n5742), .Q(n6420) );
  MUX21X1 U5516 ( .IN1(N2996), .IN2(N4121), .S(n5758), .Q(n6421) );
  MUX21X1 U5517 ( .IN1(n6421), .IN2(n5723), .S(n5742), .Q(n6422) );
  MUX41X1 U5518 ( .IN1(n6422), .IN3(n6419), .IN2(n6420), .IN4(n4444), .S0(
        n5793), .S1(n5747), .Q(n6423) );
  MUX21X1 U5519 ( .IN1(N1746), .IN2(n527), .S(n5758), .Q(n6424) );
  MUX21X1 U5520 ( .IN1(N4492), .IN2(N4525), .S(n5758), .Q(n6425) );
  MUX21X1 U5521 ( .IN1(N1779), .IN2(N1811), .S(n5757), .Q(n6426) );
  MUX41X1 U5522 ( .IN1(n6413), .IN3(n6424), .IN2(n6426), .IN4(n6425), .S0(
        n5752), .S1(n5726), .Q(n6427) );
  MUX21X1 U5523 ( .IN1(n6428), .IN2(n6427), .S(n5791), .Q(n6430) );
  MUX41X1 U5524 ( .IN1(N1811), .IN3(N1746), .IN2(N4722), .IN4(N4755), .S0(
        n5743), .S1(n5754), .Q(n6431) );
  MUX21X1 U5525 ( .IN1(n6425), .IN2(N4567), .S(n5743), .Q(n6432) );
  MUX21X1 U5526 ( .IN1(N4891), .IN2(N4959), .S(n5757), .Q(n6433) );
  AND2X1 U5527 ( .IN1(N4992), .IN2(n5778), .Q(n6434) );
  MUX21X1 U5528 ( .IN1(n6433), .IN2(n6434), .S(n5743), .Q(n6435) );
  MUX21X1 U5529 ( .IN1(n527), .IN2(N1746), .S(n5743), .Q(n6436) );
  MUX21X1 U5530 ( .IN1(n414), .IN2(n6436), .S(n5757), .Q(n6437) );
  MUX41X1 U5531 ( .IN1(n6437), .IN3(n6432), .IN2(n6435), .IN4(n6431), .S0(
        n5793), .S1(n5747), .Q(n6438) );
  MUX41X1 U5532 ( .IN1(n6438), .IN3(n6430), .IN2(n6423), .IN4(n6417), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5633) );
  MUX21X1 U5533 ( .IN1(N4785), .IN2(N4854), .S(n5757), .Q(n6439) );
  MUX21X1 U5534 ( .IN1(N1743), .IN2(n6439), .S(n5743), .Q(n6440) );
  MUX21X1 U5535 ( .IN1(N4587), .IN2(N1743), .S(n5758), .Q(n6441) );
  MUX21X1 U5536 ( .IN1(n530), .IN2(N1743), .S(n5757), .Q(n6442) );
  AND2X1 U5537 ( .IN1(N4374), .IN2(n5786), .Q(n6443) );
  MUX41X1 U5538 ( .IN1(n6443), .IN3(N5268), .IN2(n6442), .IN4(n6441), .S0(
        n5752), .S1(n5725), .Q(n6444) );
  MUX21X1 U5539 ( .IN1(n6444), .IN2(n6440), .S(n5791), .Q(n6445) );
  MUX21X1 U5540 ( .IN1(N4719), .IN2(N4752), .S(n5743), .Q(n6446) );
  MUX21X1 U5541 ( .IN1(n6446), .IN2(N1743), .S(n5757), .Q(n6447) );
  MUX21X1 U5542 ( .IN1(n530), .IN2(N5203), .S(n5743), .Q(n6448) );
  MUX21X1 U5543 ( .IN1(N2993), .IN2(N4118), .S(n5757), .Q(n6449) );
  MUX21X1 U5544 ( .IN1(n6449), .IN2(ID_imm_offset[7]), .S(n5743), .Q(n6450) );
  MUX41X1 U5545 ( .IN1(n6450), .IN3(n6447), .IN2(n6448), .IN4(n4447), .S0(
        n5793), .S1(n5747), .Q(n6451) );
  MUX21X1 U5546 ( .IN1(N1743), .IN2(n530), .S(n5757), .Q(n6452) );
  MUX21X1 U5547 ( .IN1(N4489), .IN2(N4522), .S(n5758), .Q(n6453) );
  MUX21X1 U5548 ( .IN1(N1776), .IN2(N1808), .S(n5757), .Q(n6454) );
  MUX41X1 U5549 ( .IN1(n6441), .IN3(n6452), .IN2(n6454), .IN4(n6453), .S0(
        n5752), .S1(n5724), .Q(n6455) );
  MUX21X1 U5550 ( .IN1(n6456), .IN2(n6455), .S(n5790), .Q(n6458) );
  MUX41X1 U5551 ( .IN1(N1808), .IN3(N1743), .IN2(N4719), .IN4(N4752), .S0(
        n5744), .S1(n5754), .Q(n6459) );
  MUX21X1 U5552 ( .IN1(n6453), .IN2(N4570), .S(n5742), .Q(n6460) );
  MUX21X1 U5553 ( .IN1(N4888), .IN2(N4956), .S(n5757), .Q(n6461) );
  AND2X1 U5554 ( .IN1(N4989), .IN2(n5779), .Q(n6462) );
  MUX21X1 U5555 ( .IN1(n6461), .IN2(n6462), .S(n5742), .Q(n6463) );
  MUX21X1 U5556 ( .IN1(n530), .IN2(N1743), .S(n5743), .Q(n6464) );
  MUX21X1 U5557 ( .IN1(n417), .IN2(n6464), .S(n5757), .Q(n6465) );
  MUX41X1 U5558 ( .IN1(n6465), .IN3(n6460), .IN2(n6463), .IN4(n6459), .S0(
        n5793), .S1(n5747), .Q(n6466) );
  MUX41X1 U5559 ( .IN1(n6466), .IN3(n6458), .IN2(n6451), .IN4(n6445), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5630) );
  MUX21X1 U5560 ( .IN1(N4778), .IN2(N4847), .S(n5757), .Q(n6467) );
  MUX21X1 U5561 ( .IN1(N1736), .IN2(n6467), .S(n5743), .Q(n6468) );
  MUX21X1 U5562 ( .IN1(N4580), .IN2(N1736), .S(n5757), .Q(n6469) );
  MUX21X1 U5563 ( .IN1(n537), .IN2(N1736), .S(n5756), .Q(n6470) );
  AND2X1 U5564 ( .IN1(N4381), .IN2(n5786), .Q(n6471) );
  MUX41X1 U5565 ( .IN1(n6471), .IN3(N5261), .IN2(n6470), .IN4(n6469), .S0(
        n5752), .S1(n5725), .Q(n6472) );
  MUX21X1 U5566 ( .IN1(n6472), .IN2(n6468), .S(n5790), .Q(n6473) );
  MUX21X1 U5567 ( .IN1(N4712), .IN2(N4745), .S(n5743), .Q(n6474) );
  MUX21X1 U5568 ( .IN1(n6474), .IN2(N1736), .S(n5756), .Q(n6475) );
  MUX21X1 U5569 ( .IN1(n537), .IN2(N5196), .S(n5743), .Q(n6476) );
  MUX21X1 U5570 ( .IN1(N2986), .IN2(N4111), .S(n5756), .Q(n6477) );
  MUX21X1 U5571 ( .IN1(n6477), .IN2(ID_imm_offset[0]), .S(n5743), .Q(n6478) );
  MUX41X1 U5572 ( .IN1(n6478), .IN3(n6475), .IN2(n6476), .IN4(N1254), .S0(
        n5792), .S1(n5747), .Q(n6479) );
  MUX21X1 U5573 ( .IN1(N1736), .IN2(n537), .S(n5761), .Q(n6480) );
  MUX21X1 U5574 ( .IN1(N4482), .IN2(N4515), .S(n5761), .Q(n6481) );
  MUX41X1 U5575 ( .IN1(n6469), .IN3(n6480), .IN2(n5711), .IN4(n6481), .S0(
        n5752), .S1(n5726), .Q(n6482) );
  MUX21X1 U5576 ( .IN1(n6483), .IN2(n6482), .S(n5791), .Q(n6485) );
  MUX41X1 U5577 ( .IN1(N1801), .IN3(N1736), .IN2(N4712), .IN4(N4745), .S0(
        n5695), .S1(n5754), .Q(n6486) );
  MUX21X1 U5578 ( .IN1(n6481), .IN2(N4577), .S(n5743), .Q(n6487) );
  MUX41X1 U5579 ( .IN1(N4881), .IN3(N4949), .IN2(ID_imm_offset[1]), .IN4(N4982), .S0(n5777), .S1(n5726), .Q(n6488) );
  MUX21X1 U5580 ( .IN1(n537), .IN2(N1736), .S(n5740), .Q(n6489) );
  MUX21X1 U5581 ( .IN1(n424), .IN2(n6489), .S(n5761), .Q(n6490) );
  MUX41X1 U5582 ( .IN1(n6490), .IN3(n6487), .IN2(n6488), .IN4(n6486), .S0(
        n5793), .S1(n5747), .Q(n6491) );
  MUX41X1 U5583 ( .IN1(n6491), .IN3(n6485), .IN2(n6479), .IN4(n6473), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5623) );
  MUX21X1 U5584 ( .IN1(N4779), .IN2(N4848), .S(n5761), .Q(n6492) );
  MUX21X1 U5585 ( .IN1(N1737), .IN2(n6492), .S(n5740), .Q(n6493) );
  MUX21X1 U5586 ( .IN1(N4581), .IN2(N1737), .S(n5761), .Q(n6494) );
  MUX21X1 U5587 ( .IN1(n536), .IN2(N1737), .S(n5761), .Q(n6495) );
  AND2X1 U5588 ( .IN1(N4380), .IN2(n5785), .Q(n6496) );
  MUX41X1 U5589 ( .IN1(n6496), .IN3(N5262), .IN2(n6495), .IN4(n6494), .S0(
        n5752), .S1(n5726), .Q(n6497) );
  MUX21X1 U5590 ( .IN1(n6497), .IN2(n6493), .S(n5790), .Q(n6498) );
  MUX21X1 U5591 ( .IN1(N4713), .IN2(N4746), .S(n5740), .Q(n6499) );
  MUX21X1 U5592 ( .IN1(n6499), .IN2(N1737), .S(n5761), .Q(n6500) );
  MUX21X1 U5593 ( .IN1(n536), .IN2(N5197), .S(n5740), .Q(n6501) );
  MUX21X1 U5594 ( .IN1(N2987), .IN2(N4112), .S(n5761), .Q(n6502) );
  MUX21X1 U5595 ( .IN1(n6502), .IN2(ID_imm_offset[1]), .S(n5740), .Q(n6503) );
  MUX41X1 U5596 ( .IN1(n6503), .IN3(n6500), .IN2(n6501), .IN4(n4453), .S0(
        n5792), .S1(n5746), .Q(n6504) );
  MUX21X1 U5597 ( .IN1(N1737), .IN2(n536), .S(n5761), .Q(n6505) );
  MUX21X1 U5598 ( .IN1(N4483), .IN2(N4516), .S(n5761), .Q(n6506) );
  MUX21X1 U5599 ( .IN1(N1770), .IN2(N1802), .S(n5762), .Q(n6507) );
  MUX41X1 U5600 ( .IN1(n6494), .IN3(n6505), .IN2(n6507), .IN4(n6506), .S0(
        n5752), .S1(n5728), .Q(n6508) );
  MUX21X1 U5601 ( .IN1(n6509), .IN2(n6508), .S(n5790), .Q(n6511) );
  MUX41X1 U5602 ( .IN1(N1802), .IN3(N1737), .IN2(N4713), .IN4(N4746), .S0(
        n5744), .S1(n5755), .Q(n6512) );
  MUX21X1 U5603 ( .IN1(n6506), .IN2(N4576), .S(n5740), .Q(n6513) );
  MUX41X1 U5604 ( .IN1(N4882), .IN3(N4950), .IN2(ID_imm_offset[2]), .IN4(N4983), .S0(n5777), .S1(n5727), .Q(n6514) );
  MUX21X1 U5605 ( .IN1(n536), .IN2(N1737), .S(n5740), .Q(n6515) );
  MUX21X1 U5606 ( .IN1(n423), .IN2(n6515), .S(n5762), .Q(n6516) );
  MUX41X1 U5607 ( .IN1(n6516), .IN3(n6513), .IN2(n6514), .IN4(n6512), .S0(
        n5793), .S1(n5746), .Q(n6517) );
  MUX41X1 U5608 ( .IN1(n6517), .IN3(n6511), .IN2(n6504), .IN4(n6498), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5624) );
  MUX21X1 U5609 ( .IN1(N4780), .IN2(N4849), .S(n5762), .Q(n6518) );
  MUX21X1 U5610 ( .IN1(N1738), .IN2(n6518), .S(n5740), .Q(n6519) );
  MUX21X1 U5611 ( .IN1(N4582), .IN2(N1738), .S(n5762), .Q(n6520) );
  MUX21X1 U5612 ( .IN1(n535), .IN2(N1738), .S(n5762), .Q(n6521) );
  AND2X1 U5613 ( .IN1(N4379), .IN2(n5785), .Q(n6522) );
  MUX41X1 U5614 ( .IN1(n6522), .IN3(N5263), .IN2(n6521), .IN4(n6520), .S0(
        n5752), .S1(n5728), .Q(n6523) );
  MUX21X1 U5615 ( .IN1(n6523), .IN2(n6519), .S(n5790), .Q(n6524) );
  MUX21X1 U5616 ( .IN1(N4714), .IN2(N4747), .S(n5740), .Q(n6525) );
  MUX21X1 U5617 ( .IN1(n6525), .IN2(N1738), .S(n5762), .Q(n6526) );
  MUX21X1 U5618 ( .IN1(n535), .IN2(N5198), .S(n5740), .Q(n6527) );
  MUX21X1 U5619 ( .IN1(N2988), .IN2(N4113), .S(n5762), .Q(n6528) );
  MUX21X1 U5620 ( .IN1(n6528), .IN2(ID_imm_offset[2]), .S(n5739), .Q(n6529) );
  MUX41X1 U5621 ( .IN1(n6529), .IN3(n6526), .IN2(n6527), .IN4(n4452), .S0(
        n5793), .S1(n5746), .Q(n6530) );
  MUX21X1 U5622 ( .IN1(N1738), .IN2(n535), .S(n5762), .Q(n6531) );
  MUX21X1 U5623 ( .IN1(N4484), .IN2(N4517), .S(n5762), .Q(n6532) );
  MUX21X1 U5624 ( .IN1(N1771), .IN2(N1803), .S(n5762), .Q(n6533) );
  MUX41X1 U5625 ( .IN1(n6520), .IN3(n6531), .IN2(n6533), .IN4(n6532), .S0(
        n5752), .S1(n5728), .Q(n6534) );
  MUX21X1 U5626 ( .IN1(n6535), .IN2(n6534), .S(n5789), .Q(n6537) );
  MUX41X1 U5627 ( .IN1(N1803), .IN3(N1738), .IN2(N4714), .IN4(N4747), .S0(
        n5744), .S1(n5755), .Q(n6538) );
  MUX21X1 U5628 ( .IN1(n6532), .IN2(N4575), .S(n5739), .Q(n6539) );
  MUX41X1 U5629 ( .IN1(N4883), .IN3(N4951), .IN2(ID_imm_offset[3]), .IN4(N4984), .S0(n5777), .S1(n5728), .Q(n6540) );
  MUX21X1 U5630 ( .IN1(n535), .IN2(N1738), .S(n5739), .Q(n6541) );
  MUX21X1 U5631 ( .IN1(n422), .IN2(n6541), .S(n5762), .Q(n6542) );
  MUX41X1 U5632 ( .IN1(n6542), .IN3(n6539), .IN2(n6540), .IN4(n6538), .S0(
        n5792), .S1(n5746), .Q(n6543) );
  MUX41X1 U5633 ( .IN1(n6543), .IN3(n6537), .IN2(n6530), .IN4(n6524), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5625) );
  MUX21X1 U5634 ( .IN1(N4781), .IN2(N4850), .S(n5762), .Q(n6544) );
  MUX21X1 U5635 ( .IN1(N1739), .IN2(n6544), .S(n5739), .Q(n6545) );
  MUX21X1 U5636 ( .IN1(N4583), .IN2(N1739), .S(n5762), .Q(n6546) );
  MUX21X1 U5637 ( .IN1(n534), .IN2(N1739), .S(n5762), .Q(n6547) );
  AND2X1 U5638 ( .IN1(N4378), .IN2(n5785), .Q(n6548) );
  MUX41X1 U5639 ( .IN1(n6548), .IN3(N5264), .IN2(n6547), .IN4(n6546), .S0(
        n5752), .S1(n5728), .Q(n6549) );
  MUX21X1 U5640 ( .IN1(n6549), .IN2(n6545), .S(n5789), .Q(n6550) );
  MUX21X1 U5641 ( .IN1(N4715), .IN2(N4748), .S(n5739), .Q(n6551) );
  MUX21X1 U5642 ( .IN1(n6551), .IN2(N1739), .S(n5762), .Q(n6552) );
  MUX21X1 U5643 ( .IN1(n534), .IN2(N5199), .S(n5739), .Q(n6553) );
  MUX21X1 U5644 ( .IN1(N2989), .IN2(N4114), .S(n5762), .Q(n6554) );
  MUX21X1 U5645 ( .IN1(n6554), .IN2(ID_imm_offset[3]), .S(n5739), .Q(n6555) );
  MUX41X1 U5646 ( .IN1(n6555), .IN3(n6552), .IN2(n6553), .IN4(n4451), .S0(
        n5792), .S1(n5746), .Q(n6556) );
  MUX21X1 U5647 ( .IN1(N1739), .IN2(n534), .S(n5762), .Q(n6557) );
  MUX21X1 U5648 ( .IN1(N4485), .IN2(N4518), .S(n5762), .Q(n6558) );
  MUX21X1 U5649 ( .IN1(N1772), .IN2(N1804), .S(n5763), .Q(n6559) );
  MUX41X1 U5650 ( .IN1(n6546), .IN3(n6557), .IN2(n6559), .IN4(n6558), .S0(
        n5752), .S1(n5729), .Q(n6560) );
  MUX21X1 U5651 ( .IN1(n6561), .IN2(n6560), .S(n5788), .Q(n6563) );
  MUX41X1 U5652 ( .IN1(N1804), .IN3(N1739), .IN2(N4715), .IN4(N4748), .S0(
        n5744), .S1(n5754), .Q(n6564) );
  MUX21X1 U5653 ( .IN1(n6558), .IN2(N4574), .S(n5739), .Q(n6565) );
  MUX41X1 U5654 ( .IN1(N4884), .IN3(N4952), .IN2(ID_imm_offset[4]), .IN4(N4985), .S0(n5777), .S1(n5729), .Q(n6566) );
  MUX21X1 U5655 ( .IN1(n534), .IN2(N1739), .S(n5739), .Q(n6567) );
  MUX21X1 U5656 ( .IN1(n421), .IN2(n6567), .S(n5763), .Q(n6568) );
  MUX41X1 U5657 ( .IN1(n6568), .IN3(n6565), .IN2(n6566), .IN4(n6564), .S0(
        n5793), .S1(n5746), .Q(n6569) );
  MUX41X1 U5658 ( .IN1(n6569), .IN3(n6563), .IN2(n6556), .IN4(n6550), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5626) );
  MUX21X1 U5659 ( .IN1(N4782), .IN2(N4851), .S(n5763), .Q(n6570) );
  MUX21X1 U5660 ( .IN1(N1740), .IN2(n6570), .S(n5739), .Q(n6571) );
  MUX21X1 U5661 ( .IN1(N4584), .IN2(N1740), .S(n5763), .Q(n6572) );
  MUX21X1 U5662 ( .IN1(n533), .IN2(N1740), .S(n5763), .Q(n6573) );
  AND2X1 U5663 ( .IN1(N4377), .IN2(n5782), .Q(n6574) );
  MUX41X1 U5664 ( .IN1(n6574), .IN3(N5265), .IN2(n6573), .IN4(n6572), .S0(
        n5752), .S1(n5729), .Q(n6575) );
  MUX21X1 U5665 ( .IN1(n6575), .IN2(n6571), .S(n5789), .Q(n6576) );
  MUX21X1 U5666 ( .IN1(N4716), .IN2(N4749), .S(n5739), .Q(n6577) );
  MUX21X1 U5667 ( .IN1(n6577), .IN2(N1740), .S(n5763), .Q(n6578) );
  MUX21X1 U5668 ( .IN1(n533), .IN2(N5200), .S(n5739), .Q(n6579) );
  MUX21X1 U5669 ( .IN1(N2990), .IN2(N4115), .S(n5763), .Q(n6580) );
  MUX21X1 U5670 ( .IN1(n6580), .IN2(ID_imm_offset[4]), .S(n5739), .Q(n6581) );
  MUX41X1 U5671 ( .IN1(n6581), .IN3(n6578), .IN2(n6579), .IN4(n4450), .S0(
        n5792), .S1(n5746), .Q(n6582) );
  MUX21X1 U5672 ( .IN1(N1740), .IN2(n533), .S(n5763), .Q(n6583) );
  MUX21X1 U5673 ( .IN1(N4486), .IN2(N4519), .S(n5763), .Q(n6584) );
  MUX21X1 U5674 ( .IN1(N1773), .IN2(N1805), .S(n5763), .Q(n6585) );
  MUX41X1 U5675 ( .IN1(n6572), .IN3(n6583), .IN2(n6585), .IN4(n6584), .S0(
        n5753), .S1(n5729), .Q(n6586) );
  MUX21X1 U5676 ( .IN1(n6587), .IN2(n6586), .S(n5788), .Q(n6589) );
  MUX41X1 U5677 ( .IN1(N1805), .IN3(N1740), .IN2(N4716), .IN4(N4749), .S0(
        n5744), .S1(n5755), .Q(n6590) );
  MUX21X1 U5678 ( .IN1(n6584), .IN2(N4573), .S(n5739), .Q(n6591) );
  MUX41X1 U5679 ( .IN1(N4885), .IN3(N4953), .IN2(ID_imm_offset[5]), .IN4(N4986), .S0(n5776), .S1(n5729), .Q(n6592) );
  MUX21X1 U5680 ( .IN1(n533), .IN2(N1740), .S(n5739), .Q(n6593) );
  MUX21X1 U5681 ( .IN1(n420), .IN2(n6593), .S(n5763), .Q(n6594) );
  MUX41X1 U5682 ( .IN1(n6594), .IN3(n6591), .IN2(n6592), .IN4(n6590), .S0(
        n5792), .S1(n5745), .Q(n6595) );
  MUX41X1 U5683 ( .IN1(n6595), .IN3(n6589), .IN2(n6582), .IN4(n6576), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5627) );
  MUX21X1 U5684 ( .IN1(N4783), .IN2(N4852), .S(n5763), .Q(n6596) );
  MUX21X1 U5685 ( .IN1(N1741), .IN2(n6596), .S(n5739), .Q(n6597) );
  MUX21X1 U5686 ( .IN1(N4585), .IN2(N1741), .S(n5763), .Q(n6598) );
  MUX21X1 U5687 ( .IN1(n532), .IN2(N1741), .S(n5763), .Q(n6599) );
  AND2X1 U5688 ( .IN1(N4376), .IN2(n5784), .Q(n6600) );
  MUX41X1 U5689 ( .IN1(n6600), .IN3(N5266), .IN2(n6599), .IN4(n6598), .S0(
        n5753), .S1(n5728), .Q(n6601) );
  MUX21X1 U5690 ( .IN1(n6601), .IN2(n6597), .S(n5788), .Q(n6602) );
  MUX21X1 U5691 ( .IN1(N4717), .IN2(N4750), .S(n5739), .Q(n6603) );
  MUX21X1 U5692 ( .IN1(n6603), .IN2(N1741), .S(n5763), .Q(n6604) );
  MUX21X1 U5693 ( .IN1(n532), .IN2(N5201), .S(n5739), .Q(n6605) );
  MUX21X1 U5694 ( .IN1(N2991), .IN2(N4116), .S(n5763), .Q(n6606) );
  MUX21X1 U5695 ( .IN1(n6606), .IN2(ID_imm_offset[5]), .S(n5738), .Q(n6607) );
  MUX41X1 U5696 ( .IN1(n6607), .IN3(n6604), .IN2(n6605), .IN4(n4449), .S0(
        n5793), .S1(n5745), .Q(n6608) );
  MUX21X1 U5697 ( .IN1(N1741), .IN2(n532), .S(n5763), .Q(n6609) );
  MUX21X1 U5698 ( .IN1(N4487), .IN2(N4520), .S(n5763), .Q(n6610) );
  MUX21X1 U5699 ( .IN1(N1774), .IN2(N1806), .S(n5764), .Q(n6611) );
  MUX41X1 U5700 ( .IN1(n6598), .IN3(n6609), .IN2(n6611), .IN4(n6610), .S0(
        n5753), .S1(n5727), .Q(n6612) );
  MUX21X1 U5701 ( .IN1(n6613), .IN2(n6612), .S(n5788), .Q(n6615) );
  MUX41X1 U5702 ( .IN1(N1806), .IN3(N1741), .IN2(N4717), .IN4(N4750), .S0(
        n5744), .S1(n5756), .Q(n6616) );
  MUX21X1 U5703 ( .IN1(n6610), .IN2(N4572), .S(n5738), .Q(n6617) );
  MUX41X1 U5704 ( .IN1(N4886), .IN3(N4954), .IN2(ID_imm_offset[6]), .IN4(N4987), .S0(n5777), .S1(n5727), .Q(n6618) );
  MUX21X1 U5705 ( .IN1(n532), .IN2(N1741), .S(n5738), .Q(n6619) );
  MUX21X1 U5706 ( .IN1(n419), .IN2(n6619), .S(n5764), .Q(n6620) );
  MUX41X1 U5707 ( .IN1(n6620), .IN3(n6617), .IN2(n6618), .IN4(n6616), .S0(
        n5792), .S1(n5745), .Q(n6621) );
  MUX41X1 U5708 ( .IN1(n6621), .IN3(n6615), .IN2(n6608), .IN4(n6602), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5628) );
  MUX21X1 U5709 ( .IN1(N4784), .IN2(N4853), .S(n5764), .Q(n6622) );
  MUX21X1 U5710 ( .IN1(N1742), .IN2(n6622), .S(n5738), .Q(n6623) );
  MUX21X1 U5711 ( .IN1(N4586), .IN2(N1742), .S(n5764), .Q(n6624) );
  MUX21X1 U5712 ( .IN1(n531), .IN2(N1742), .S(n5764), .Q(n6625) );
  AND2X1 U5713 ( .IN1(N4375), .IN2(n5783), .Q(n6626) );
  MUX41X1 U5714 ( .IN1(n6626), .IN3(N5267), .IN2(n6625), .IN4(n6624), .S0(
        n5753), .S1(n5726), .Q(n6627) );
  MUX21X1 U5715 ( .IN1(n6627), .IN2(n6623), .S(n5787), .Q(n6628) );
  MUX21X1 U5716 ( .IN1(N4718), .IN2(N4751), .S(n5738), .Q(n6629) );
  MUX21X1 U5717 ( .IN1(n6629), .IN2(N1742), .S(n5764), .Q(n6630) );
  MUX21X1 U5718 ( .IN1(n531), .IN2(N5202), .S(n5738), .Q(n6631) );
  MUX21X1 U5719 ( .IN1(N2992), .IN2(N4117), .S(n5764), .Q(n6632) );
  MUX21X1 U5720 ( .IN1(n6632), .IN2(ID_imm_offset[6]), .S(n5738), .Q(n6633) );
  MUX41X1 U5721 ( .IN1(n6633), .IN3(n6630), .IN2(n6631), .IN4(n4448), .S0(
        n5792), .S1(n5745), .Q(n6634) );
  MUX21X1 U5722 ( .IN1(N1742), .IN2(n531), .S(n5764), .Q(n6635) );
  MUX21X1 U5723 ( .IN1(N4488), .IN2(N4521), .S(n5764), .Q(n6636) );
  MUX21X1 U5724 ( .IN1(N1775), .IN2(N1807), .S(n5764), .Q(n6637) );
  MUX41X1 U5725 ( .IN1(n6624), .IN3(n6635), .IN2(n6637), .IN4(n6636), .S0(
        n5752), .S1(n5727), .Q(n6638) );
  MUX21X1 U5726 ( .IN1(n6639), .IN2(n6638), .S(n5787), .Q(n6641) );
  MUX41X1 U5727 ( .IN1(N1807), .IN3(N1742), .IN2(N4718), .IN4(N4751), .S0(
        n5744), .S1(n5755), .Q(n6642) );
  MUX21X1 U5728 ( .IN1(n6636), .IN2(N4571), .S(n5738), .Q(n6643) );
  MUX41X1 U5729 ( .IN1(N4887), .IN3(N4955), .IN2(ID_imm_offset[7]), .IN4(N4988), .S0(n5776), .S1(n5727), .Q(n6644) );
  MUX21X1 U5730 ( .IN1(n531), .IN2(N1742), .S(n5738), .Q(n6645) );
  MUX21X1 U5731 ( .IN1(n418), .IN2(n6645), .S(n5764), .Q(n6646) );
  MUX41X1 U5732 ( .IN1(n6646), .IN3(n6643), .IN2(n6644), .IN4(n6642), .S0(
        n5793), .S1(n5745), .Q(n6647) );
  MUX41X1 U5733 ( .IN1(n6647), .IN3(n6641), .IN2(n6634), .IN4(n6628), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5629) );
  MUX21X1 U5734 ( .IN1(N4777), .IN2(N4846), .S(n5764), .Q(n6648) );
  MUX21X1 U5735 ( .IN1(N1735), .IN2(n6648), .S(n5738), .Q(n6649) );
  MUX21X1 U5736 ( .IN1(N4579), .IN2(N1735), .S(n5764), .Q(n6650) );
  MUX21X1 U5737 ( .IN1(n538), .IN2(N1735), .S(n5764), .Q(n6651) );
  AND2X1 U5738 ( .IN1(N4382), .IN2(n5781), .Q(n6652) );
  MUX41X1 U5739 ( .IN1(n6652), .IN3(N5260), .IN2(n6651), .IN4(n6650), .S0(
        n5753), .S1(n5727), .Q(n6653) );
  MUX21X1 U5740 ( .IN1(n6653), .IN2(n6649), .S(n5787), .Q(n6654) );
  MUX21X1 U5741 ( .IN1(N4711), .IN2(N4744), .S(n5738), .Q(n6655) );
  MUX21X1 U5742 ( .IN1(n6655), .IN2(N1735), .S(n5764), .Q(n6656) );
  MUX21X1 U5743 ( .IN1(n538), .IN2(N5195), .S(n5738), .Q(n6657) );
  AND2X1 U5744 ( .IN1(n6659), .IN2(n3723), .Q(n6658) );
  MUX41X1 U5745 ( .IN1(n6658), .IN3(n6656), .IN2(n6657), .IN4(N1255), .S0(
        n5792), .S1(n5745), .Q(n6660) );
  MUX21X1 U5746 ( .IN1(N1735), .IN2(n538), .S(n5764), .Q(n6661) );
  MUX21X1 U5747 ( .IN1(N4481), .IN2(N4514), .S(n5764), .Q(n6662) );
  MUX41X1 U5748 ( .IN1(n6650), .IN3(n6661), .IN2(n5712), .IN4(n6662), .S0(
        n5752), .S1(n5725), .Q(n6663) );
  MUX21X1 U5749 ( .IN1(n6664), .IN2(n6663), .S(n5787), .Q(n6666) );
  MUX41X1 U5750 ( .IN1(N1800), .IN3(N1735), .IN2(N4711), .IN4(N4744), .S0(
        n5744), .S1(n5754), .Q(n6667) );
  MUX21X1 U5751 ( .IN1(n6662), .IN2(N4578), .S(n5738), .Q(n6668) );
  MUX41X1 U5752 ( .IN1(N4880), .IN3(N4948), .IN2(ID_imm_offset[0]), .IN4(N4981), .S0(n5777), .S1(n5726), .Q(n6669) );
  MUX21X1 U5753 ( .IN1(n538), .IN2(N1735), .S(n5738), .Q(n6670) );
  MUX21X1 U5754 ( .IN1(n425), .IN2(n6670), .S(n5764), .Q(n6671) );
  MUX41X1 U5755 ( .IN1(n6671), .IN3(n6668), .IN2(n6669), .IN4(n6667), .S0(
        n5793), .S1(n5745), .Q(n6672) );
  MUX41X1 U5756 ( .IN1(n6672), .IN3(n6666), .IN2(n6660), .IN4(n6654), .S0(
        ID_opcode[2]), .S1(ID_opcode[3]), .Q(N5622) );
  OR2X1 U5757 ( .IN1(N5055), .IN2(n5777), .Q(n6673) );
  OR2X1 U5758 ( .IN1(N5054), .IN2(n5777), .Q(n6674) );
  OR2X1 U5759 ( .IN1(N5053), .IN2(n5777), .Q(n6675) );
  OR2X1 U5760 ( .IN1(N5052), .IN2(n5777), .Q(n6676) );
  OR2X1 U5761 ( .IN1(N5051), .IN2(n5777), .Q(n6677) );
  OR2X1 U5762 ( .IN1(N5050), .IN2(n5777), .Q(n6678) );
  OR2X1 U5763 ( .IN1(N5049), .IN2(n5777), .Q(n6679) );
  OR2X1 U5764 ( .IN1(N5048), .IN2(n5777), .Q(n6680) );
  OR2X1 U5765 ( .IN1(N5047), .IN2(n5777), .Q(n6681) );
  OR2X1 U5766 ( .IN1(N5046), .IN2(n5777), .Q(n6682) );
  OR2X1 U5767 ( .IN1(N5058), .IN2(n5777), .Q(n6683) );
  OR2X1 U5768 ( .IN1(N5065), .IN2(n5778), .Q(n6684) );
  OR2X1 U5769 ( .IN1(N5064), .IN2(n5777), .Q(n6685) );
  OR2X1 U5770 ( .IN1(N5063), .IN2(n5777), .Q(n6686) );
  OR2X1 U5771 ( .IN1(N5062), .IN2(n5777), .Q(n6687) );
  OR2X1 U5772 ( .IN1(N5061), .IN2(n5778), .Q(n6688) );
  OR2X1 U5773 ( .IN1(N5060), .IN2(n5777), .Q(n6689) );
  OR2X1 U5774 ( .IN1(N5059), .IN2(n5778), .Q(n6690) );
  OR2X1 U5775 ( .IN1(N5057), .IN2(n5777), .Q(n6691) );
  OR2X1 U5776 ( .IN1(N5056), .IN2(n5778), .Q(n6692) );
  OR2X1 U5777 ( .IN1(N5068), .IN2(n5778), .Q(n6693) );
  OR2X1 U5778 ( .IN1(N5067), .IN2(n5778), .Q(n6694) );
  OR2X1 U5779 ( .IN1(N5066), .IN2(n5778), .Q(n6695) );
  OR2X1 U5780 ( .IN1(N5069), .IN2(n5778), .Q(n6696) );
  OR2X1 U5781 ( .IN1(N5076), .IN2(n5778), .Q(n6697) );
  OR2X1 U5782 ( .IN1(N5075), .IN2(n5778), .Q(n6698) );
  OR2X1 U5783 ( .IN1(N5074), .IN2(n5778), .Q(n6699) );
  OR2X1 U5784 ( .IN1(N5073), .IN2(n5778), .Q(n6700) );
  OR2X1 U5785 ( .IN1(N5072), .IN2(n5778), .Q(n6701) );
  OR2X1 U5786 ( .IN1(N5071), .IN2(n5778), .Q(n6702) );
  OR2X1 U5787 ( .IN1(N5070), .IN2(n5778), .Q(n6703) );
  OR2X1 U5788 ( .IN1(N5077), .IN2(n5778), .Q(n6704) );
  MUX21X1 U5789 ( .IN1(n4463), .IN2(n403), .S(n5765), .Q(n6705) );
  MUX21X1 U5790 ( .IN1(n6705), .IN2(n6673), .S(n5738), .Q(n5815) );
  MUX21X1 U5791 ( .IN1(n4462), .IN2(n402), .S(n5765), .Q(n6706) );
  MUX21X1 U5792 ( .IN1(n6706), .IN2(n6674), .S(n5738), .Q(n5843) );
  MUX21X1 U5793 ( .IN1(n4461), .IN2(n401), .S(n5765), .Q(n6707) );
  MUX21X1 U5794 ( .IN1(n6707), .IN2(n6675), .S(n5738), .Q(n5871) );
  MUX21X1 U5795 ( .IN1(n4460), .IN2(n400), .S(n5765), .Q(n6708) );
  MUX21X1 U5796 ( .IN1(n6708), .IN2(n6676), .S(n5738), .Q(n5899) );
  MUX21X1 U5797 ( .IN1(n4459), .IN2(n399), .S(n5765), .Q(n6709) );
  MUX21X1 U5798 ( .IN1(n6709), .IN2(n6677), .S(n5737), .Q(n5927) );
  MUX21X1 U5799 ( .IN1(n4458), .IN2(n398), .S(n5765), .Q(n6710) );
  MUX21X1 U5800 ( .IN1(n6710), .IN2(n6678), .S(n5737), .Q(n5955) );
  MUX21X1 U5801 ( .IN1(n4457), .IN2(n397), .S(n5765), .Q(n6711) );
  MUX21X1 U5802 ( .IN1(n6711), .IN2(n6679), .S(n5737), .Q(n5983) );
  MUX21X1 U5803 ( .IN1(n4456), .IN2(n396), .S(n5765), .Q(n6712) );
  MUX21X1 U5804 ( .IN1(n6712), .IN2(n6680), .S(n5737), .Q(n6011) );
  MUX21X1 U5805 ( .IN1(n4455), .IN2(n395), .S(n5765), .Q(n6713) );
  MUX21X1 U5806 ( .IN1(n6713), .IN2(n6681), .S(n5737), .Q(n6039) );
  MUX21X1 U5807 ( .IN1(n4454), .IN2(n394), .S(n5765), .Q(n6714) );
  MUX21X1 U5808 ( .IN1(n6714), .IN2(n6682), .S(n5737), .Q(n6067) );
  MUX21X1 U5809 ( .IN1(n4466), .IN2(n406), .S(n5765), .Q(n6715) );
  MUX21X1 U5810 ( .IN1(n6715), .IN2(n6683), .S(n5737), .Q(n6095) );
  MUX21X1 U5811 ( .IN1(n4473), .IN2(n413), .S(n5765), .Q(n6716) );
  MUX21X1 U5812 ( .IN1(n6716), .IN2(n6684), .S(n5737), .Q(n6123) );
  MUX21X1 U5813 ( .IN1(n4472), .IN2(n412), .S(n5765), .Q(n6717) );
  MUX21X1 U5814 ( .IN1(n6717), .IN2(n6685), .S(n5737), .Q(n6151) );
  MUX21X1 U5815 ( .IN1(n4471), .IN2(n411), .S(n5765), .Q(n6718) );
  MUX21X1 U5816 ( .IN1(n6718), .IN2(n6686), .S(n5737), .Q(n6179) );
  MUX21X1 U5817 ( .IN1(n4470), .IN2(n410), .S(n5765), .Q(n6719) );
  MUX21X1 U5818 ( .IN1(n6719), .IN2(n6687), .S(n5737), .Q(n6207) );
  MUX21X1 U5819 ( .IN1(n4469), .IN2(n409), .S(n5765), .Q(n6720) );
  MUX21X1 U5820 ( .IN1(n6720), .IN2(n6688), .S(n5737), .Q(n6235) );
  MUX21X1 U5821 ( .IN1(n4468), .IN2(n408), .S(n5765), .Q(n6721) );
  MUX21X1 U5822 ( .IN1(n6721), .IN2(n6689), .S(n5737), .Q(n6263) );
  MUX21X1 U5823 ( .IN1(n4467), .IN2(n407), .S(n5766), .Q(n6722) );
  MUX21X1 U5824 ( .IN1(n6722), .IN2(n6690), .S(n5737), .Q(n6291) );
  MUX21X1 U5825 ( .IN1(n4465), .IN2(n405), .S(n5766), .Q(n6723) );
  MUX21X1 U5826 ( .IN1(n6723), .IN2(n6691), .S(n5737), .Q(n6319) );
  MUX21X1 U5827 ( .IN1(n4464), .IN2(n404), .S(n5766), .Q(n6724) );
  MUX21X1 U5828 ( .IN1(n6724), .IN2(n6692), .S(n5737), .Q(n6347) );
  MUX21X1 U5829 ( .IN1(n4476), .IN2(n416), .S(n5766), .Q(n6725) );
  MUX21X1 U5830 ( .IN1(n6725), .IN2(n6693), .S(n5737), .Q(n6374) );
  MUX21X1 U5831 ( .IN1(n4475), .IN2(n415), .S(n5766), .Q(n6726) );
  MUX21X1 U5832 ( .IN1(n6726), .IN2(n6694), .S(n5737), .Q(n6401) );
  MUX21X1 U5833 ( .IN1(n4474), .IN2(n414), .S(n5766), .Q(n6727) );
  MUX21X1 U5834 ( .IN1(n6727), .IN2(n6695), .S(n5736), .Q(n6429) );
  MUX21X1 U5835 ( .IN1(n4477), .IN2(n417), .S(n5766), .Q(n6728) );
  MUX21X1 U5836 ( .IN1(n6728), .IN2(n6696), .S(n5736), .Q(n6457) );
  MUX21X1 U5837 ( .IN1(n4484), .IN2(n424), .S(n5766), .Q(n6729) );
  MUX21X1 U5838 ( .IN1(n6729), .IN2(n6697), .S(n5736), .Q(n6484) );
  MUX21X1 U5839 ( .IN1(n4483), .IN2(n423), .S(n5766), .Q(n6730) );
  MUX21X1 U5840 ( .IN1(n6730), .IN2(n6698), .S(n5736), .Q(n6510) );
  MUX21X1 U5841 ( .IN1(n4482), .IN2(n422), .S(n5766), .Q(n6731) );
  MUX21X1 U5842 ( .IN1(n6731), .IN2(n6699), .S(n5736), .Q(n6536) );
  MUX21X1 U5843 ( .IN1(n4481), .IN2(n421), .S(n5766), .Q(n6732) );
  MUX21X1 U5844 ( .IN1(n6732), .IN2(n6700), .S(n5736), .Q(n6562) );
  MUX21X1 U5845 ( .IN1(n4480), .IN2(n420), .S(n5766), .Q(n6733) );
  MUX21X1 U5846 ( .IN1(n6733), .IN2(n6701), .S(n5736), .Q(n6588) );
  MUX21X1 U5847 ( .IN1(n4479), .IN2(n419), .S(n5766), .Q(n6734) );
  MUX21X1 U5848 ( .IN1(n6734), .IN2(n6702), .S(n5736), .Q(n6614) );
  MUX21X1 U5849 ( .IN1(n4478), .IN2(n418), .S(n5766), .Q(n6735) );
  MUX21X1 U5850 ( .IN1(n6735), .IN2(n6703), .S(n5740), .Q(n6640) );
  MUX21X1 U5851 ( .IN1(N2985), .IN2(N4110), .S(n5766), .Q(n6659) );
  MUX21X1 U5852 ( .IN1(n4485), .IN2(n425), .S(n5766), .Q(n6736) );
  MUX21X1 U5853 ( .IN1(n6736), .IN2(n6704), .S(n5730), .Q(n6665) );
  MUX41X1 U5854 ( .IN1(\R[4][0] ), .IN3(\R[6][0] ), .IN2(\R[5][0] ), .IN4(
        \R[7][0] ), .S0(N307), .S1(n6801), .Q(n6737) );
  MUX41X1 U5855 ( .IN1(\R[0][0] ), .IN3(\R[2][0] ), .IN2(\R[1][0] ), .IN4(
        \R[3][0] ), .S0(N307), .S1(n6807), .Q(n6738) );
  MUX21X1 U5856 ( .IN1(n6738), .IN2(n6737), .S(N308), .Q(N498) );
  MUX41X1 U5857 ( .IN1(\R[4][1] ), .IN3(\R[6][1] ), .IN2(\R[5][1] ), .IN4(
        \R[7][1] ), .S0(N307), .S1(n6804), .Q(n6739) );
  MUX41X1 U5858 ( .IN1(\R[0][1] ), .IN3(\R[2][1] ), .IN2(\R[1][1] ), .IN4(
        \R[3][1] ), .S0(N307), .S1(n6801), .Q(n6740) );
  MUX21X1 U5859 ( .IN1(n6740), .IN2(n6739), .S(N308), .Q(N497) );
  MUX41X1 U5860 ( .IN1(\R[4][2] ), .IN3(\R[6][2] ), .IN2(\R[5][2] ), .IN4(
        \R[7][2] ), .S0(N307), .S1(n6803), .Q(n6741) );
  MUX41X1 U5861 ( .IN1(\R[0][2] ), .IN3(\R[2][2] ), .IN2(\R[1][2] ), .IN4(
        \R[3][2] ), .S0(N307), .S1(n6805), .Q(n6742) );
  MUX21X1 U5862 ( .IN1(n6742), .IN2(n6741), .S(N308), .Q(N496) );
  MUX41X1 U5863 ( .IN1(\R[4][3] ), .IN3(\R[6][3] ), .IN2(\R[5][3] ), .IN4(
        \R[7][3] ), .S0(N307), .S1(n6801), .Q(n6743) );
  MUX41X1 U5864 ( .IN1(\R[0][3] ), .IN3(\R[2][3] ), .IN2(\R[1][3] ), .IN4(
        \R[3][3] ), .S0(N307), .S1(n6806), .Q(n6744) );
  MUX21X1 U5865 ( .IN1(n6744), .IN2(n6743), .S(N308), .Q(N495) );
  MUX41X1 U5866 ( .IN1(\R[4][4] ), .IN3(\R[6][4] ), .IN2(\R[5][4] ), .IN4(
        \R[7][4] ), .S0(N307), .S1(n6807), .Q(n6745) );
  MUX41X1 U5867 ( .IN1(\R[0][4] ), .IN3(\R[2][4] ), .IN2(\R[1][4] ), .IN4(
        \R[3][4] ), .S0(N307), .S1(n6807), .Q(n6746) );
  MUX21X1 U5868 ( .IN1(n6746), .IN2(n6745), .S(N308), .Q(N494) );
  MUX41X1 U5869 ( .IN1(\R[4][5] ), .IN3(\R[6][5] ), .IN2(\R[5][5] ), .IN4(
        \R[7][5] ), .S0(N307), .S1(n6806), .Q(n6747) );
  MUX41X1 U5870 ( .IN1(\R[0][5] ), .IN3(\R[2][5] ), .IN2(\R[1][5] ), .IN4(
        \R[3][5] ), .S0(N307), .S1(n6806), .Q(n6748) );
  MUX21X1 U5871 ( .IN1(n6748), .IN2(n6747), .S(N308), .Q(N493) );
  MUX41X1 U5872 ( .IN1(\R[4][6] ), .IN3(\R[6][6] ), .IN2(\R[5][6] ), .IN4(
        \R[7][6] ), .S0(N307), .S1(n6805), .Q(n6749) );
  MUX41X1 U5873 ( .IN1(\R[0][6] ), .IN3(\R[2][6] ), .IN2(\R[1][6] ), .IN4(
        \R[3][6] ), .S0(N307), .S1(n6805), .Q(n6750) );
  MUX21X1 U5874 ( .IN1(n6750), .IN2(n6749), .S(N308), .Q(N492) );
  MUX41X1 U5875 ( .IN1(\R[4][7] ), .IN3(\R[6][7] ), .IN2(\R[5][7] ), .IN4(
        \R[7][7] ), .S0(N307), .S1(n6806), .Q(n6751) );
  MUX41X1 U5876 ( .IN1(\R[0][7] ), .IN3(\R[2][7] ), .IN2(\R[1][7] ), .IN4(
        \R[3][7] ), .S0(N307), .S1(n6804), .Q(n6752) );
  MUX21X1 U5877 ( .IN1(n6752), .IN2(n6751), .S(N308), .Q(N491) );
  MUX41X1 U5878 ( .IN1(\R[4][8] ), .IN3(\R[6][8] ), .IN2(\R[5][8] ), .IN4(
        \R[7][8] ), .S0(N307), .S1(n6805), .Q(n6753) );
  MUX41X1 U5879 ( .IN1(\R[0][8] ), .IN3(\R[2][8] ), .IN2(\R[1][8] ), .IN4(
        \R[3][8] ), .S0(N307), .S1(n6803), .Q(n6754) );
  MUX21X1 U5880 ( .IN1(n6754), .IN2(n6753), .S(N308), .Q(N490) );
  MUX41X1 U5881 ( .IN1(\R[4][9] ), .IN3(\R[6][9] ), .IN2(\R[5][9] ), .IN4(
        \R[7][9] ), .S0(N307), .S1(n5699), .Q(n6755) );
  MUX41X1 U5882 ( .IN1(\R[0][9] ), .IN3(\R[2][9] ), .IN2(\R[1][9] ), .IN4(
        \R[3][9] ), .S0(N307), .S1(n6802), .Q(n6756) );
  MUX21X1 U5883 ( .IN1(n6756), .IN2(n6755), .S(N308), .Q(N489) );
  MUX41X1 U5884 ( .IN1(\R[4][10] ), .IN3(\R[6][10] ), .IN2(\R[5][10] ), .IN4(
        \R[7][10] ), .S0(N307), .S1(n5699), .Q(n6757) );
  MUX41X1 U5885 ( .IN1(\R[0][10] ), .IN3(\R[2][10] ), .IN2(\R[1][10] ), .IN4(
        \R[3][10] ), .S0(N307), .S1(n6801), .Q(n6758) );
  MUX21X1 U5886 ( .IN1(n6758), .IN2(n6757), .S(N308), .Q(N488) );
  MUX41X1 U5887 ( .IN1(\R[4][11] ), .IN3(\R[6][11] ), .IN2(\R[5][11] ), .IN4(
        \R[7][11] ), .S0(N307), .S1(n6806), .Q(n6759) );
  MUX41X1 U5888 ( .IN1(\R[0][11] ), .IN3(\R[2][11] ), .IN2(\R[1][11] ), .IN4(
        \R[3][11] ), .S0(N307), .S1(n6805), .Q(n6760) );
  MUX21X1 U5889 ( .IN1(n6760), .IN2(n6759), .S(N308), .Q(N487) );
  MUX41X1 U5890 ( .IN1(\R[4][12] ), .IN3(\R[6][12] ), .IN2(\R[5][12] ), .IN4(
        \R[7][12] ), .S0(N307), .S1(n6802), .Q(n6761) );
  MUX41X1 U5891 ( .IN1(\R[0][12] ), .IN3(\R[2][12] ), .IN2(\R[1][12] ), .IN4(
        \R[3][12] ), .S0(N307), .S1(n5699), .Q(n6762) );
  MUX21X1 U5892 ( .IN1(n6762), .IN2(n6761), .S(N308), .Q(N486) );
  MUX41X1 U5893 ( .IN1(\R[4][13] ), .IN3(\R[6][13] ), .IN2(\R[5][13] ), .IN4(
        \R[7][13] ), .S0(N307), .S1(n6804), .Q(n6763) );
  MUX41X1 U5894 ( .IN1(\R[0][13] ), .IN3(\R[2][13] ), .IN2(\R[1][13] ), .IN4(
        \R[3][13] ), .S0(N307), .S1(n6807), .Q(n6764) );
  MUX21X1 U5895 ( .IN1(n6764), .IN2(n6763), .S(N308), .Q(N485) );
  MUX41X1 U5896 ( .IN1(\R[4][14] ), .IN3(\R[6][14] ), .IN2(\R[5][14] ), .IN4(
        \R[7][14] ), .S0(N307), .S1(n6801), .Q(n6765) );
  MUX41X1 U5897 ( .IN1(\R[0][14] ), .IN3(\R[2][14] ), .IN2(\R[1][14] ), .IN4(
        \R[3][14] ), .S0(N307), .S1(n6802), .Q(n6766) );
  MUX21X1 U5898 ( .IN1(n6766), .IN2(n6765), .S(N308), .Q(N484) );
  MUX41X1 U5899 ( .IN1(\R[4][15] ), .IN3(\R[6][15] ), .IN2(\R[5][15] ), .IN4(
        \R[7][15] ), .S0(N307), .S1(n6805), .Q(n6767) );
  MUX21X1 U5900 ( .IN1(n6768), .IN2(n6767), .S(N308), .Q(N483) );
  MUX41X1 U5901 ( .IN1(\R[4][16] ), .IN3(\R[6][16] ), .IN2(\R[5][16] ), .IN4(
        \R[7][16] ), .S0(N307), .S1(n6803), .Q(n6769) );
  MUX41X1 U5902 ( .IN1(\R[0][16] ), .IN3(\R[2][16] ), .IN2(\R[1][16] ), .IN4(
        \R[3][16] ), .S0(N307), .S1(n5699), .Q(n6770) );
  MUX21X1 U5903 ( .IN1(n6770), .IN2(n6769), .S(N308), .Q(N482) );
  MUX41X1 U5904 ( .IN1(\R[4][17] ), .IN3(\R[6][17] ), .IN2(\R[5][17] ), .IN4(
        \R[7][17] ), .S0(N307), .S1(n6801), .Q(n6771) );
  MUX21X1 U5905 ( .IN1(n6772), .IN2(n6771), .S(N308), .Q(N481) );
  MUX41X1 U5906 ( .IN1(\R[4][18] ), .IN3(\R[6][18] ), .IN2(\R[5][18] ), .IN4(
        \R[7][18] ), .S0(N307), .S1(n6802), .Q(n6773) );
  MUX41X1 U5907 ( .IN1(\R[0][18] ), .IN3(\R[2][18] ), .IN2(\R[1][18] ), .IN4(
        \R[3][18] ), .S0(N307), .S1(n6803), .Q(n6774) );
  MUX21X1 U5908 ( .IN1(n6774), .IN2(n6773), .S(N308), .Q(N480) );
  MUX41X1 U5909 ( .IN1(\R[4][19] ), .IN3(\R[6][19] ), .IN2(\R[5][19] ), .IN4(
        \R[7][19] ), .S0(N307), .S1(n5699), .Q(n6775) );
  MUX21X1 U5910 ( .IN1(n6776), .IN2(n6775), .S(N308), .Q(N479) );
  MUX41X1 U5911 ( .IN1(\R[4][20] ), .IN3(\R[6][20] ), .IN2(\R[5][20] ), .IN4(
        \R[7][20] ), .S0(N307), .S1(n6804), .Q(n6777) );
  MUX41X1 U5912 ( .IN1(\R[0][20] ), .IN3(\R[2][20] ), .IN2(\R[1][20] ), .IN4(
        \R[3][20] ), .S0(N307), .S1(n6807), .Q(n6778) );
  MUX21X1 U5913 ( .IN1(n6778), .IN2(n6777), .S(N308), .Q(N478) );
  MUX41X1 U5914 ( .IN1(\R[4][21] ), .IN3(\R[6][21] ), .IN2(\R[5][21] ), .IN4(
        \R[7][21] ), .S0(N307), .S1(n6805), .Q(n6779) );
  MUX21X1 U5915 ( .IN1(n6780), .IN2(n6779), .S(N308), .Q(N477) );
  MUX41X1 U5916 ( .IN1(\R[4][22] ), .IN3(\R[6][22] ), .IN2(\R[5][22] ), .IN4(
        \R[7][22] ), .S0(N307), .S1(n5699), .Q(n6781) );
  MUX41X1 U5917 ( .IN1(\R[0][22] ), .IN3(\R[2][22] ), .IN2(\R[1][22] ), .IN4(
        \R[3][22] ), .S0(N307), .S1(n6804), .Q(n6782) );
  MUX21X1 U5918 ( .IN1(n6782), .IN2(n6781), .S(N308), .Q(N476) );
  MUX41X1 U5919 ( .IN1(\R[4][23] ), .IN3(\R[6][23] ), .IN2(\R[5][23] ), .IN4(
        \R[7][23] ), .S0(N307), .S1(n6803), .Q(n6783) );
  MUX21X1 U5920 ( .IN1(n6784), .IN2(n6783), .S(N308), .Q(N475) );
  MUX41X1 U5921 ( .IN1(\R[4][24] ), .IN3(\R[6][24] ), .IN2(\R[5][24] ), .IN4(
        \R[7][24] ), .S0(N307), .S1(n6806), .Q(n6785) );
  MUX41X1 U5922 ( .IN1(\R[0][24] ), .IN3(\R[2][24] ), .IN2(\R[1][24] ), .IN4(
        \R[3][24] ), .S0(N307), .S1(n6806), .Q(n6786) );
  MUX21X1 U5923 ( .IN1(n6786), .IN2(n6785), .S(N308), .Q(N474) );
  MUX41X1 U5924 ( .IN1(\R[4][25] ), .IN3(\R[6][25] ), .IN2(\R[5][25] ), .IN4(
        \R[7][25] ), .S0(N307), .S1(n6807), .Q(n6787) );
  MUX41X1 U5925 ( .IN1(\R[0][25] ), .IN3(\R[2][25] ), .IN2(\R[1][25] ), .IN4(
        \R[3][25] ), .S0(N307), .S1(n6802), .Q(n6788) );
  MUX21X1 U5926 ( .IN1(n6788), .IN2(n6787), .S(N308), .Q(N473) );
  MUX41X1 U5927 ( .IN1(\R[4][26] ), .IN3(\R[6][26] ), .IN2(\R[5][26] ), .IN4(
        \R[7][26] ), .S0(N307), .S1(n6807), .Q(n6789) );
  MUX21X1 U5928 ( .IN1(n6790), .IN2(n6789), .S(N308), .Q(N472) );
  MUX41X1 U5929 ( .IN1(\R[4][27] ), .IN3(\R[6][27] ), .IN2(\R[5][27] ), .IN4(
        \R[7][27] ), .S0(N307), .S1(n6804), .Q(n6791) );
  MUX41X1 U5930 ( .IN1(\R[0][27] ), .IN3(\R[2][27] ), .IN2(\R[1][27] ), .IN4(
        \R[3][27] ), .S0(N307), .S1(n6802), .Q(n6792) );
  MUX21X1 U5931 ( .IN1(n6792), .IN2(n6791), .S(N308), .Q(N471) );
  MUX41X1 U5932 ( .IN1(\R[4][28] ), .IN3(\R[6][28] ), .IN2(\R[5][28] ), .IN4(
        \R[7][28] ), .S0(N307), .S1(n6803), .Q(n6793) );
  MUX21X1 U5933 ( .IN1(n6794), .IN2(n6793), .S(N308), .Q(N470) );
  MUX41X1 U5934 ( .IN1(\R[4][29] ), .IN3(\R[6][29] ), .IN2(\R[5][29] ), .IN4(
        \R[7][29] ), .S0(N307), .S1(n6802), .Q(n6795) );
  MUX41X1 U5935 ( .IN1(\R[0][29] ), .IN3(\R[2][29] ), .IN2(\R[1][29] ), .IN4(
        \R[3][29] ), .S0(N307), .S1(n6801), .Q(n6796) );
  MUX21X1 U5936 ( .IN1(n6796), .IN2(n6795), .S(N308), .Q(N469) );
  MUX41X1 U5937 ( .IN1(\R[4][30] ), .IN3(\R[6][30] ), .IN2(\R[5][30] ), .IN4(
        \R[7][30] ), .S0(N307), .S1(n6804), .Q(n6797) );
  MUX21X1 U5938 ( .IN1(n6798), .IN2(n6797), .S(N308), .Q(N468) );
  MUX41X1 U5939 ( .IN1(\R[4][31] ), .IN3(\R[6][31] ), .IN2(\R[5][31] ), .IN4(
        \R[7][31] ), .S0(N307), .S1(n6803), .Q(n6799) );
  MUX41X1 U5940 ( .IN1(\R[0][31] ), .IN3(\R[2][31] ), .IN2(\R[1][31] ), .IN4(
        \R[3][31] ), .S0(N307), .S1(n5699), .Q(n6800) );
  MUX21X1 U5941 ( .IN1(n6800), .IN2(n6799), .S(N308), .Q(N467) );
  MUX41X1 U5942 ( .IN1(\R[4][0] ), .IN3(\R[6][0] ), .IN2(\R[5][0] ), .IN4(
        \R[7][0] ), .S0(N310), .S1(n6874), .Q(n6808) );
  MUX41X1 U5943 ( .IN1(\R[0][0] ), .IN3(\R[2][0] ), .IN2(\R[1][0] ), .IN4(
        \R[3][0] ), .S0(N310), .S1(n6875), .Q(n6809) );
  MUX21X1 U5944 ( .IN1(n6809), .IN2(n6808), .S(N311), .Q(N530) );
  MUX41X1 U5945 ( .IN1(\R[4][1] ), .IN3(\R[6][1] ), .IN2(\R[5][1] ), .IN4(
        \R[7][1] ), .S0(N310), .S1(n6876), .Q(n6810) );
  MUX21X1 U5946 ( .IN1(n6811), .IN2(n6810), .S(N311), .Q(N529) );
  MUX41X1 U5947 ( .IN1(\R[4][2] ), .IN3(\R[6][2] ), .IN2(\R[5][2] ), .IN4(
        \R[7][2] ), .S0(N310), .S1(n6874), .Q(n6812) );
  MUX41X1 U5948 ( .IN1(\R[0][2] ), .IN3(\R[2][2] ), .IN2(\R[1][2] ), .IN4(
        \R[3][2] ), .S0(N310), .S1(n6874), .Q(n6813) );
  MUX21X1 U5949 ( .IN1(n6813), .IN2(n6812), .S(N311), .Q(N528) );
  MUX41X1 U5950 ( .IN1(\R[4][3] ), .IN3(\R[6][3] ), .IN2(\R[5][3] ), .IN4(
        \R[7][3] ), .S0(N310), .S1(n7333), .Q(n6814) );
  MUX21X1 U5951 ( .IN1(n6815), .IN2(n6814), .S(N311), .Q(N527) );
  MUX41X1 U5952 ( .IN1(\R[4][4] ), .IN3(\R[6][4] ), .IN2(\R[5][4] ), .IN4(
        \R[7][4] ), .S0(N310), .S1(n7333), .Q(n6816) );
  MUX41X1 U5953 ( .IN1(\R[0][4] ), .IN3(\R[2][4] ), .IN2(\R[1][4] ), .IN4(
        \R[3][4] ), .S0(N310), .S1(n6877), .Q(n6817) );
  MUX21X1 U5954 ( .IN1(n6817), .IN2(n6816), .S(N311), .Q(N526) );
  MUX41X1 U5955 ( .IN1(\R[4][5] ), .IN3(\R[6][5] ), .IN2(\R[5][5] ), .IN4(
        \R[7][5] ), .S0(N310), .S1(n6872), .Q(n6818) );
  MUX21X1 U5956 ( .IN1(n6819), .IN2(n6818), .S(N311), .Q(N525) );
  MUX41X1 U5957 ( .IN1(\R[4][6] ), .IN3(\R[6][6] ), .IN2(\R[5][6] ), .IN4(
        \R[7][6] ), .S0(N310), .S1(n6872), .Q(n6820) );
  MUX41X1 U5958 ( .IN1(\R[0][6] ), .IN3(\R[2][6] ), .IN2(\R[1][6] ), .IN4(
        \R[3][6] ), .S0(N310), .S1(n7333), .Q(n6821) );
  MUX21X1 U5959 ( .IN1(n6821), .IN2(n6820), .S(N311), .Q(N524) );
  MUX41X1 U5960 ( .IN1(\R[4][7] ), .IN3(\R[6][7] ), .IN2(\R[5][7] ), .IN4(
        \R[7][7] ), .S0(N310), .S1(n6873), .Q(n6822) );
  MUX41X1 U5961 ( .IN1(\R[0][7] ), .IN3(\R[2][7] ), .IN2(\R[1][7] ), .IN4(
        \R[3][7] ), .S0(N310), .S1(n6873), .Q(n6823) );
  MUX21X1 U5962 ( .IN1(n6823), .IN2(n6822), .S(N311), .Q(N523) );
  MUX41X1 U5963 ( .IN1(\R[4][8] ), .IN3(\R[6][8] ), .IN2(\R[5][8] ), .IN4(
        \R[7][8] ), .S0(N310), .S1(n6874), .Q(n6824) );
  MUX21X1 U5964 ( .IN1(n6825), .IN2(n6824), .S(N311), .Q(N522) );
  MUX41X1 U5965 ( .IN1(\R[4][9] ), .IN3(\R[6][9] ), .IN2(\R[5][9] ), .IN4(
        \R[7][9] ), .S0(N310), .S1(n5698), .Q(n6826) );
  MUX41X1 U5966 ( .IN1(\R[0][9] ), .IN3(\R[2][9] ), .IN2(\R[1][9] ), .IN4(
        \R[3][9] ), .S0(N310), .S1(n6873), .Q(n6827) );
  MUX21X1 U5967 ( .IN1(n6827), .IN2(n6826), .S(N311), .Q(N521) );
  MUX41X1 U5968 ( .IN1(\R[4][10] ), .IN3(\R[6][10] ), .IN2(\R[5][10] ), .IN4(
        \R[7][10] ), .S0(N310), .S1(n6877), .Q(n6828) );
  MUX21X1 U5969 ( .IN1(n6829), .IN2(n6828), .S(N311), .Q(N520) );
  MUX41X1 U5970 ( .IN1(\R[4][11] ), .IN3(\R[6][11] ), .IN2(\R[5][11] ), .IN4(
        \R[7][11] ), .S0(N310), .S1(n6875), .Q(n6830) );
  MUX41X1 U5971 ( .IN1(\R[0][11] ), .IN3(\R[2][11] ), .IN2(\R[1][11] ), .IN4(
        \R[3][11] ), .S0(N310), .S1(n6877), .Q(n6831) );
  MUX21X1 U5972 ( .IN1(n6831), .IN2(n6830), .S(N311), .Q(N519) );
  MUX41X1 U5973 ( .IN1(\R[4][12] ), .IN3(\R[6][12] ), .IN2(\R[5][12] ), .IN4(
        \R[7][12] ), .S0(N310), .S1(n6877), .Q(n6832) );
  MUX21X1 U5974 ( .IN1(n6833), .IN2(n6832), .S(N311), .Q(N518) );
  MUX41X1 U5975 ( .IN1(\R[4][13] ), .IN3(\R[6][13] ), .IN2(\R[5][13] ), .IN4(
        \R[7][13] ), .S0(N310), .S1(n7333), .Q(n6834) );
  MUX41X1 U5976 ( .IN1(\R[0][13] ), .IN3(\R[2][13] ), .IN2(\R[1][13] ), .IN4(
        \R[3][13] ), .S0(N310), .S1(n6876), .Q(n6835) );
  MUX21X1 U5977 ( .IN1(n6835), .IN2(n6834), .S(N311), .Q(N517) );
  MUX41X1 U5978 ( .IN1(\R[4][14] ), .IN3(\R[6][14] ), .IN2(\R[5][14] ), .IN4(
        \R[7][14] ), .S0(N310), .S1(n6876), .Q(n6836) );
  MUX21X1 U5979 ( .IN1(n6837), .IN2(n6836), .S(N311), .Q(N516) );
  MUX41X1 U5980 ( .IN1(\R[4][15] ), .IN3(\R[6][15] ), .IN2(\R[5][15] ), .IN4(
        \R[7][15] ), .S0(N310), .S1(n6872), .Q(n6838) );
  MUX41X1 U5981 ( .IN1(\R[0][15] ), .IN3(\R[2][15] ), .IN2(\R[1][15] ), .IN4(
        \R[3][15] ), .S0(N310), .S1(n6875), .Q(n6839) );
  MUX21X1 U5982 ( .IN1(n6839), .IN2(n6838), .S(N311), .Q(N515) );
  MUX41X1 U5983 ( .IN1(\R[4][16] ), .IN3(\R[6][16] ), .IN2(\R[5][16] ), .IN4(
        \R[7][16] ), .S0(N310), .S1(n6876), .Q(n6840) );
  MUX21X1 U5984 ( .IN1(n6841), .IN2(n6840), .S(N311), .Q(N514) );
  MUX41X1 U5985 ( .IN1(\R[4][17] ), .IN3(\R[6][17] ), .IN2(\R[5][17] ), .IN4(
        \R[7][17] ), .S0(N310), .S1(n6877), .Q(n6842) );
  MUX41X1 U5986 ( .IN1(\R[0][17] ), .IN3(\R[2][17] ), .IN2(\R[1][17] ), .IN4(
        \R[3][17] ), .S0(N310), .S1(n6874), .Q(n6843) );
  MUX21X1 U5987 ( .IN1(n6843), .IN2(n6842), .S(N311), .Q(N513) );
  MUX41X1 U5988 ( .IN1(\R[4][18] ), .IN3(\R[6][18] ), .IN2(\R[5][18] ), .IN4(
        \R[7][18] ), .S0(N310), .S1(n6872), .Q(n6844) );
  MUX41X1 U5989 ( .IN1(\R[0][18] ), .IN3(\R[2][18] ), .IN2(\R[1][18] ), .IN4(
        \R[3][18] ), .S0(N310), .S1(n6873), .Q(n6845) );
  MUX21X1 U5990 ( .IN1(n6845), .IN2(n6844), .S(N311), .Q(N512) );
  MUX41X1 U5991 ( .IN1(\R[4][19] ), .IN3(\R[6][19] ), .IN2(\R[5][19] ), .IN4(
        \R[7][19] ), .S0(N310), .S1(n6872), .Q(n6846) );
  MUX41X1 U5992 ( .IN1(\R[0][19] ), .IN3(\R[2][19] ), .IN2(\R[1][19] ), .IN4(
        \R[3][19] ), .S0(N310), .S1(n6872), .Q(n6847) );
  MUX21X1 U5993 ( .IN1(n6847), .IN2(n6846), .S(N311), .Q(N511) );
  MUX41X1 U5994 ( .IN1(\R[4][20] ), .IN3(\R[6][20] ), .IN2(\R[5][20] ), .IN4(
        \R[7][20] ), .S0(N310), .S1(n6873), .Q(n6848) );
  MUX41X1 U5995 ( .IN1(\R[0][20] ), .IN3(\R[2][20] ), .IN2(\R[1][20] ), .IN4(
        \R[3][20] ), .S0(N310), .S1(n5698), .Q(n6849) );
  MUX21X1 U5996 ( .IN1(n6849), .IN2(n6848), .S(N311), .Q(N510) );
  MUX41X1 U5997 ( .IN1(\R[4][21] ), .IN3(\R[6][21] ), .IN2(\R[5][21] ), .IN4(
        \R[7][21] ), .S0(N310), .S1(n5698), .Q(n6850) );
  MUX41X1 U5998 ( .IN1(\R[0][21] ), .IN3(\R[2][21] ), .IN2(\R[1][21] ), .IN4(
        \R[3][21] ), .S0(N310), .S1(n6877), .Q(n6851) );
  MUX21X1 U5999 ( .IN1(n6851), .IN2(n6850), .S(N311), .Q(N509) );
  MUX41X1 U6000 ( .IN1(\R[4][22] ), .IN3(\R[6][22] ), .IN2(\R[5][22] ), .IN4(
        \R[7][22] ), .S0(N310), .S1(n7333), .Q(n6852) );
  MUX41X1 U6001 ( .IN1(\R[0][22] ), .IN3(\R[2][22] ), .IN2(\R[1][22] ), .IN4(
        \R[3][22] ), .S0(N310), .S1(n6873), .Q(n6853) );
  MUX21X1 U6002 ( .IN1(n6853), .IN2(n6852), .S(N311), .Q(N508) );
  MUX41X1 U6003 ( .IN1(\R[4][23] ), .IN3(\R[6][23] ), .IN2(\R[5][23] ), .IN4(
        \R[7][23] ), .S0(N310), .S1(n6877), .Q(n6854) );
  MUX41X1 U6004 ( .IN1(\R[0][23] ), .IN3(\R[2][23] ), .IN2(\R[1][23] ), .IN4(
        \R[3][23] ), .S0(N310), .S1(n5698), .Q(n6855) );
  MUX21X1 U6005 ( .IN1(n6855), .IN2(n6854), .S(N311), .Q(N507) );
  MUX41X1 U6006 ( .IN1(\R[4][24] ), .IN3(\R[6][24] ), .IN2(\R[5][24] ), .IN4(
        \R[7][24] ), .S0(N310), .S1(n6876), .Q(n6856) );
  MUX41X1 U6007 ( .IN1(\R[0][24] ), .IN3(\R[2][24] ), .IN2(\R[1][24] ), .IN4(
        \R[3][24] ), .S0(N310), .S1(n6873), .Q(n6857) );
  MUX21X1 U6008 ( .IN1(n6857), .IN2(n6856), .S(N311), .Q(N506) );
  MUX41X1 U6009 ( .IN1(\R[4][25] ), .IN3(\R[6][25] ), .IN2(\R[5][25] ), .IN4(
        \R[7][25] ), .S0(N310), .S1(n6876), .Q(n6858) );
  MUX41X1 U6010 ( .IN1(\R[0][25] ), .IN3(\R[2][25] ), .IN2(\R[1][25] ), .IN4(
        \R[3][25] ), .S0(N310), .S1(n6875), .Q(n6859) );
  MUX21X1 U6011 ( .IN1(n6859), .IN2(n6858), .S(N311), .Q(N505) );
  MUX41X1 U6012 ( .IN1(\R[4][26] ), .IN3(\R[6][26] ), .IN2(\R[5][26] ), .IN4(
        \R[7][26] ), .S0(N310), .S1(n6874), .Q(n6860) );
  MUX41X1 U6013 ( .IN1(\R[0][26] ), .IN3(\R[2][26] ), .IN2(\R[1][26] ), .IN4(
        \R[3][26] ), .S0(N310), .S1(n7333), .Q(n6861) );
  MUX21X1 U6014 ( .IN1(n6861), .IN2(n6860), .S(N311), .Q(N504) );
  MUX41X1 U6015 ( .IN1(\R[4][27] ), .IN3(\R[6][27] ), .IN2(\R[5][27] ), .IN4(
        \R[7][27] ), .S0(N310), .S1(n6874), .Q(n6862) );
  MUX41X1 U6016 ( .IN1(\R[0][27] ), .IN3(\R[2][27] ), .IN2(\R[1][27] ), .IN4(
        \R[3][27] ), .S0(N310), .S1(n6875), .Q(n6863) );
  MUX21X1 U6017 ( .IN1(n6863), .IN2(n6862), .S(N311), .Q(N503) );
  MUX41X1 U6018 ( .IN1(\R[4][28] ), .IN3(\R[6][28] ), .IN2(\R[5][28] ), .IN4(
        \R[7][28] ), .S0(N310), .S1(n6872), .Q(n6864) );
  MUX41X1 U6019 ( .IN1(\R[0][28] ), .IN3(\R[2][28] ), .IN2(\R[1][28] ), .IN4(
        \R[3][28] ), .S0(N310), .S1(n6876), .Q(n6865) );
  MUX21X1 U6020 ( .IN1(n6865), .IN2(n6864), .S(N311), .Q(N502) );
  MUX41X1 U6021 ( .IN1(\R[4][29] ), .IN3(\R[6][29] ), .IN2(\R[5][29] ), .IN4(
        \R[7][29] ), .S0(N310), .S1(n5698), .Q(n6866) );
  MUX41X1 U6022 ( .IN1(\R[0][29] ), .IN3(\R[2][29] ), .IN2(\R[1][29] ), .IN4(
        \R[3][29] ), .S0(N310), .S1(n6875), .Q(n6867) );
  MUX21X1 U6023 ( .IN1(n6867), .IN2(n6866), .S(N311), .Q(N501) );
  MUX41X1 U6024 ( .IN1(\R[4][30] ), .IN3(\R[6][30] ), .IN2(\R[5][30] ), .IN4(
        \R[7][30] ), .S0(N310), .S1(n6877), .Q(n6868) );
  MUX41X1 U6025 ( .IN1(\R[0][30] ), .IN3(\R[2][30] ), .IN2(\R[1][30] ), .IN4(
        \R[3][30] ), .S0(N310), .S1(n6875), .Q(n6869) );
  MUX21X1 U6026 ( .IN1(n6869), .IN2(n6868), .S(N311), .Q(N500) );
  MUX41X1 U6027 ( .IN1(\R[4][31] ), .IN3(\R[6][31] ), .IN2(\R[5][31] ), .IN4(
        \R[7][31] ), .S0(N310), .S1(n5698), .Q(n6870) );
  MUX41X1 U6028 ( .IN1(\R[0][31] ), .IN3(\R[2][31] ), .IN2(\R[1][31] ), .IN4(
        \R[3][31] ), .S0(N310), .S1(n5698), .Q(n6871) );
  MUX21X1 U6029 ( .IN1(n6871), .IN2(n6870), .S(N311), .Q(N499) );
  MUX41X1 U6030 ( .IN1(\R[4][0] ), .IN3(\R[6][0] ), .IN2(\R[5][0] ), .IN4(
        \R[7][0] ), .S0(N313), .S1(n6950), .Q(n6878) );
  MUX41X1 U6031 ( .IN1(\R[0][0] ), .IN3(\R[2][0] ), .IN2(\R[1][0] ), .IN4(
        \R[3][0] ), .S0(N313), .S1(n6949), .Q(n6879) );
  MUX21X1 U6032 ( .IN1(n6879), .IN2(n6878), .S(n7022), .Q(N562) );
  MUX41X1 U6033 ( .IN1(\R[4][1] ), .IN3(\R[6][1] ), .IN2(\R[5][1] ), .IN4(
        \R[7][1] ), .S0(N313), .S1(n6948), .Q(n6880) );
  MUX41X1 U6034 ( .IN1(\R[0][1] ), .IN3(\R[2][1] ), .IN2(\R[1][1] ), .IN4(
        \R[3][1] ), .S0(N313), .S1(n6947), .Q(n6881) );
  MUX21X1 U6035 ( .IN1(n6881), .IN2(n6880), .S(n7019), .Q(N561) );
  MUX41X1 U6036 ( .IN1(\R[4][2] ), .IN3(\R[6][2] ), .IN2(\R[5][2] ), .IN4(
        \R[7][2] ), .S0(N313), .S1(n6946), .Q(n6882) );
  MUX41X1 U6037 ( .IN1(\R[0][2] ), .IN3(\R[2][2] ), .IN2(\R[1][2] ), .IN4(
        \R[3][2] ), .S0(N313), .S1(n6945), .Q(n6883) );
  MUX21X1 U6038 ( .IN1(n6883), .IN2(n6882), .S(n7016), .Q(N560) );
  MUX41X1 U6039 ( .IN1(\R[4][3] ), .IN3(\R[6][3] ), .IN2(\R[5][3] ), .IN4(
        \R[7][3] ), .S0(N313), .S1(n6944), .Q(n6884) );
  MUX41X1 U6040 ( .IN1(\R[0][3] ), .IN3(\R[2][3] ), .IN2(\R[1][3] ), .IN4(
        \R[3][3] ), .S0(N313), .S1(n6943), .Q(n6885) );
  MUX21X1 U6041 ( .IN1(n6885), .IN2(n6884), .S(n7015), .Q(N559) );
  MUX41X1 U6042 ( .IN1(\R[4][4] ), .IN3(\R[6][4] ), .IN2(\R[5][4] ), .IN4(
        \R[7][4] ), .S0(N313), .S1(n6943), .Q(n6886) );
  MUX41X1 U6043 ( .IN1(\R[0][4] ), .IN3(\R[2][4] ), .IN2(\R[1][4] ), .IN4(
        \R[3][4] ), .S0(N313), .S1(n6942), .Q(n6887) );
  MUX21X1 U6044 ( .IN1(n6887), .IN2(n6886), .S(n7021), .Q(N558) );
  MUX41X1 U6045 ( .IN1(\R[4][5] ), .IN3(\R[6][5] ), .IN2(\R[5][5] ), .IN4(
        \R[7][5] ), .S0(N313), .S1(n5700), .Q(n6888) );
  MUX41X1 U6046 ( .IN1(\R[0][5] ), .IN3(\R[2][5] ), .IN2(\R[1][5] ), .IN4(
        \R[3][5] ), .S0(N313), .S1(n6948), .Q(n6889) );
  MUX21X1 U6047 ( .IN1(n6889), .IN2(n6888), .S(n7022), .Q(N557) );
  MUX41X1 U6048 ( .IN1(\R[4][6] ), .IN3(\R[6][6] ), .IN2(\R[5][6] ), .IN4(
        \R[7][6] ), .S0(N313), .S1(n6943), .Q(n6890) );
  MUX41X1 U6049 ( .IN1(\R[0][6] ), .IN3(\R[2][6] ), .IN2(\R[1][6] ), .IN4(
        \R[3][6] ), .S0(N313), .S1(n6944), .Q(n6891) );
  MUX21X1 U6050 ( .IN1(n6891), .IN2(n6890), .S(n7024), .Q(N556) );
  MUX41X1 U6051 ( .IN1(\R[4][7] ), .IN3(\R[6][7] ), .IN2(\R[5][7] ), .IN4(
        \R[7][7] ), .S0(N313), .S1(n6950), .Q(n6892) );
  MUX41X1 U6052 ( .IN1(\R[0][7] ), .IN3(\R[2][7] ), .IN2(\R[1][7] ), .IN4(
        \R[3][7] ), .S0(N313), .S1(n6949), .Q(n6893) );
  MUX21X1 U6053 ( .IN1(n6893), .IN2(n6892), .S(n7026), .Q(N555) );
  MUX41X1 U6054 ( .IN1(\R[4][8] ), .IN3(\R[6][8] ), .IN2(\R[5][8] ), .IN4(
        \R[7][8] ), .S0(N313), .S1(n6942), .Q(n6894) );
  MUX41X1 U6055 ( .IN1(\R[0][8] ), .IN3(\R[2][8] ), .IN2(\R[1][8] ), .IN4(
        \R[3][8] ), .S0(N313), .S1(n6948), .Q(n6895) );
  MUX21X1 U6056 ( .IN1(n6895), .IN2(n6894), .S(n7017), .Q(N554) );
  MUX41X1 U6057 ( .IN1(\R[4][9] ), .IN3(\R[6][9] ), .IN2(\R[5][9] ), .IN4(
        \R[7][9] ), .S0(N313), .S1(n6947), .Q(n6896) );
  MUX41X1 U6058 ( .IN1(\R[0][9] ), .IN3(\R[2][9] ), .IN2(\R[1][9] ), .IN4(
        \R[3][9] ), .S0(N313), .S1(n6947), .Q(n6897) );
  MUX21X1 U6059 ( .IN1(n6897), .IN2(n6896), .S(n7017), .Q(N553) );
  MUX41X1 U6060 ( .IN1(\R[4][10] ), .IN3(\R[6][10] ), .IN2(\R[5][10] ), .IN4(
        \R[7][10] ), .S0(N313), .S1(n5700), .Q(n6898) );
  MUX41X1 U6061 ( .IN1(\R[0][10] ), .IN3(\R[2][10] ), .IN2(\R[1][10] ), .IN4(
        \R[3][10] ), .S0(N313), .S1(n6946), .Q(n6899) );
  MUX21X1 U6062 ( .IN1(n6899), .IN2(n6898), .S(n7020), .Q(N552) );
  MUX41X1 U6063 ( .IN1(\R[4][11] ), .IN3(\R[6][11] ), .IN2(\R[5][11] ), .IN4(
        \R[7][11] ), .S0(N313), .S1(n6944), .Q(n6900) );
  MUX41X1 U6064 ( .IN1(\R[0][11] ), .IN3(\R[2][11] ), .IN2(\R[1][11] ), .IN4(
        \R[3][11] ), .S0(N313), .S1(n6946), .Q(n6901) );
  MUX21X1 U6065 ( .IN1(n6901), .IN2(n6900), .S(n7019), .Q(N551) );
  MUX41X1 U6066 ( .IN1(\R[4][12] ), .IN3(\R[6][12] ), .IN2(\R[5][12] ), .IN4(
        \R[7][12] ), .S0(N313), .S1(n6949), .Q(n6902) );
  MUX41X1 U6067 ( .IN1(\R[0][12] ), .IN3(\R[2][12] ), .IN2(\R[1][12] ), .IN4(
        \R[3][12] ), .S0(N313), .S1(n6948), .Q(n6903) );
  MUX21X1 U6068 ( .IN1(n6903), .IN2(n6902), .S(n7025), .Q(N550) );
  MUX41X1 U6069 ( .IN1(\R[4][13] ), .IN3(\R[6][13] ), .IN2(\R[5][13] ), .IN4(
        \R[7][13] ), .S0(N313), .S1(n6942), .Q(n6904) );
  MUX41X1 U6070 ( .IN1(\R[0][13] ), .IN3(\R[2][13] ), .IN2(\R[1][13] ), .IN4(
        \R[3][13] ), .S0(N313), .S1(n5700), .Q(n6905) );
  MUX21X1 U6071 ( .IN1(n6905), .IN2(n6904), .S(n7021), .Q(N549) );
  MUX41X1 U6072 ( .IN1(\R[4][14] ), .IN3(\R[6][14] ), .IN2(\R[5][14] ), .IN4(
        \R[7][14] ), .S0(N313), .S1(n6945), .Q(n6906) );
  MUX41X1 U6073 ( .IN1(\R[0][14] ), .IN3(\R[2][14] ), .IN2(\R[1][14] ), .IN4(
        \R[3][14] ), .S0(N313), .S1(n6944), .Q(n6907) );
  MUX21X1 U6074 ( .IN1(n6907), .IN2(n6906), .S(n7022), .Q(N548) );
  MUX41X1 U6075 ( .IN1(\R[4][15] ), .IN3(\R[6][15] ), .IN2(\R[5][15] ), .IN4(
        \R[7][15] ), .S0(N313), .S1(n6943), .Q(n6908) );
  MUX41X1 U6076 ( .IN1(\R[0][15] ), .IN3(\R[2][15] ), .IN2(\R[1][15] ), .IN4(
        \R[3][15] ), .S0(N313), .S1(n6947), .Q(n6909) );
  MUX21X1 U6077 ( .IN1(n6909), .IN2(n6908), .S(n7021), .Q(N547) );
  MUX41X1 U6078 ( .IN1(\R[4][16] ), .IN3(\R[6][16] ), .IN2(\R[5][16] ), .IN4(
        \R[7][16] ), .S0(N313), .S1(n6947), .Q(n6910) );
  MUX41X1 U6079 ( .IN1(\R[0][16] ), .IN3(\R[2][16] ), .IN2(\R[1][16] ), .IN4(
        \R[3][16] ), .S0(N313), .S1(n6945), .Q(n6911) );
  MUX21X1 U6080 ( .IN1(n6911), .IN2(n6910), .S(n7024), .Q(N546) );
  MUX41X1 U6081 ( .IN1(\R[4][17] ), .IN3(\R[6][17] ), .IN2(\R[5][17] ), .IN4(
        \R[7][17] ), .S0(N313), .S1(n6949), .Q(n6912) );
  MUX41X1 U6082 ( .IN1(\R[0][17] ), .IN3(\R[2][17] ), .IN2(\R[1][17] ), .IN4(
        \R[3][17] ), .S0(N313), .S1(n6950), .Q(n6913) );
  MUX21X1 U6083 ( .IN1(n6913), .IN2(n6912), .S(n7023), .Q(N545) );
  MUX41X1 U6084 ( .IN1(\R[4][18] ), .IN3(\R[6][18] ), .IN2(\R[5][18] ), .IN4(
        \R[7][18] ), .S0(N313), .S1(n6946), .Q(n6914) );
  MUX41X1 U6085 ( .IN1(\R[0][18] ), .IN3(\R[2][18] ), .IN2(\R[1][18] ), .IN4(
        \R[3][18] ), .S0(N313), .S1(n6943), .Q(n6915) );
  MUX21X1 U6086 ( .IN1(n6915), .IN2(n6914), .S(n7026), .Q(N544) );
  MUX41X1 U6087 ( .IN1(\R[4][19] ), .IN3(\R[6][19] ), .IN2(\R[5][19] ), .IN4(
        \R[7][19] ), .S0(N313), .S1(n6942), .Q(n6916) );
  MUX41X1 U6088 ( .IN1(\R[0][19] ), .IN3(\R[2][19] ), .IN2(\R[1][19] ), .IN4(
        \R[3][19] ), .S0(N313), .S1(n5700), .Q(n6917) );
  MUX21X1 U6089 ( .IN1(n6917), .IN2(n6916), .S(n7025), .Q(N543) );
  MUX41X1 U6090 ( .IN1(\R[4][20] ), .IN3(\R[6][20] ), .IN2(\R[5][20] ), .IN4(
        \R[7][20] ), .S0(N313), .S1(n6947), .Q(n6918) );
  MUX41X1 U6091 ( .IN1(\R[0][20] ), .IN3(\R[2][20] ), .IN2(\R[1][20] ), .IN4(
        \R[3][20] ), .S0(N313), .S1(n6942), .Q(n6919) );
  MUX21X1 U6092 ( .IN1(n6919), .IN2(n6918), .S(n7021), .Q(N542) );
  MUX41X1 U6093 ( .IN1(\R[4][21] ), .IN3(\R[6][21] ), .IN2(\R[5][21] ), .IN4(
        \R[7][21] ), .S0(N313), .S1(n6946), .Q(n6920) );
  MUX41X1 U6094 ( .IN1(\R[0][21] ), .IN3(\R[2][21] ), .IN2(\R[1][21] ), .IN4(
        \R[3][21] ), .S0(N313), .S1(n6948), .Q(n6921) );
  MUX21X1 U6095 ( .IN1(n6921), .IN2(n6920), .S(n5697), .Q(N541) );
  MUX41X1 U6096 ( .IN1(\R[4][22] ), .IN3(\R[6][22] ), .IN2(\R[5][22] ), .IN4(
        \R[7][22] ), .S0(N313), .S1(n6944), .Q(n6922) );
  MUX41X1 U6097 ( .IN1(\R[0][22] ), .IN3(\R[2][22] ), .IN2(\R[1][22] ), .IN4(
        \R[3][22] ), .S0(N313), .S1(n6944), .Q(n6923) );
  MUX21X1 U6098 ( .IN1(n6923), .IN2(n6922), .S(n7024), .Q(N540) );
  MUX41X1 U6099 ( .IN1(\R[4][23] ), .IN3(\R[6][23] ), .IN2(\R[5][23] ), .IN4(
        \R[7][23] ), .S0(N313), .S1(n6944), .Q(n6924) );
  MUX41X1 U6100 ( .IN1(\R[0][23] ), .IN3(\R[2][23] ), .IN2(\R[1][23] ), .IN4(
        \R[3][23] ), .S0(N313), .S1(n6949), .Q(n6925) );
  MUX21X1 U6101 ( .IN1(n6925), .IN2(n6924), .S(n7018), .Q(N539) );
  MUX41X1 U6102 ( .IN1(\R[4][24] ), .IN3(\R[6][24] ), .IN2(\R[5][24] ), .IN4(
        \R[7][24] ), .S0(N313), .S1(n6945), .Q(n6926) );
  MUX41X1 U6103 ( .IN1(\R[0][24] ), .IN3(\R[2][24] ), .IN2(\R[1][24] ), .IN4(
        \R[3][24] ), .S0(N313), .S1(n6943), .Q(n6927) );
  MUX21X1 U6104 ( .IN1(n6927), .IN2(n6926), .S(n7018), .Q(N538) );
  MUX41X1 U6105 ( .IN1(\R[4][25] ), .IN3(\R[6][25] ), .IN2(\R[5][25] ), .IN4(
        \R[7][25] ), .S0(N313), .S1(n6945), .Q(n6928) );
  MUX41X1 U6106 ( .IN1(\R[0][25] ), .IN3(\R[2][25] ), .IN2(\R[1][25] ), .IN4(
        \R[3][25] ), .S0(N313), .S1(n6950), .Q(n6929) );
  MUX21X1 U6107 ( .IN1(n6929), .IN2(n6928), .S(n5697), .Q(N537) );
  MUX41X1 U6108 ( .IN1(\R[4][26] ), .IN3(\R[6][26] ), .IN2(\R[5][26] ), .IN4(
        \R[7][26] ), .S0(N313), .S1(n6950), .Q(n6930) );
  MUX41X1 U6109 ( .IN1(\R[0][26] ), .IN3(\R[2][26] ), .IN2(\R[1][26] ), .IN4(
        \R[3][26] ), .S0(N313), .S1(n6946), .Q(n6931) );
  MUX21X1 U6110 ( .IN1(n6931), .IN2(n6930), .S(n7021), .Q(N536) );
  MUX41X1 U6111 ( .IN1(\R[4][27] ), .IN3(\R[6][27] ), .IN2(\R[5][27] ), .IN4(
        \R[7][27] ), .S0(N313), .S1(n6942), .Q(n6932) );
  MUX41X1 U6112 ( .IN1(\R[0][27] ), .IN3(\R[2][27] ), .IN2(\R[1][27] ), .IN4(
        \R[3][27] ), .S0(N313), .S1(n6948), .Q(n6933) );
  MUX21X1 U6113 ( .IN1(n6933), .IN2(n6932), .S(n7018), .Q(N535) );
  MUX41X1 U6114 ( .IN1(\R[4][28] ), .IN3(\R[6][28] ), .IN2(\R[5][28] ), .IN4(
        \R[7][28] ), .S0(N313), .S1(n6943), .Q(n6934) );
  MUX41X1 U6115 ( .IN1(\R[0][28] ), .IN3(\R[2][28] ), .IN2(\R[1][28] ), .IN4(
        \R[3][28] ), .S0(N313), .S1(n5700), .Q(n6935) );
  MUX21X1 U6116 ( .IN1(n6935), .IN2(n6934), .S(n7026), .Q(N534) );
  MUX41X1 U6117 ( .IN1(\R[4][29] ), .IN3(\R[6][29] ), .IN2(\R[5][29] ), .IN4(
        \R[7][29] ), .S0(N313), .S1(n6945), .Q(n6936) );
  MUX41X1 U6118 ( .IN1(\R[0][29] ), .IN3(\R[2][29] ), .IN2(\R[1][29] ), .IN4(
        \R[3][29] ), .S0(N313), .S1(n6942), .Q(n6937) );
  MUX21X1 U6119 ( .IN1(n6937), .IN2(n6936), .S(n5697), .Q(N533) );
  MUX41X1 U6120 ( .IN1(\R[4][30] ), .IN3(\R[6][30] ), .IN2(\R[5][30] ), .IN4(
        \R[7][30] ), .S0(N313), .S1(n6950), .Q(n6938) );
  MUX41X1 U6121 ( .IN1(\R[0][30] ), .IN3(\R[2][30] ), .IN2(\R[1][30] ), .IN4(
        \R[3][30] ), .S0(N313), .S1(n6949), .Q(n6939) );
  MUX21X1 U6122 ( .IN1(n6939), .IN2(n6938), .S(n5697), .Q(N532) );
  MUX41X1 U6123 ( .IN1(\R[4][31] ), .IN3(\R[6][31] ), .IN2(\R[5][31] ), .IN4(
        \R[7][31] ), .S0(N313), .S1(n5700), .Q(n6940) );
  MUX41X1 U6124 ( .IN1(\R[0][31] ), .IN3(\R[2][31] ), .IN2(\R[1][31] ), .IN4(
        \R[3][31] ), .S0(N313), .S1(n5700), .Q(n6941) );
  MUX21X1 U6125 ( .IN1(n6941), .IN2(n6940), .S(n5697), .Q(N531) );
  MUX41X1 U6126 ( .IN1(\R[4][0] ), .IN3(\R[6][0] ), .IN2(\R[5][0] ), .IN4(
        \R[7][0] ), .S0(N136), .S1(n7023), .Q(n6951) );
  MUX41X1 U6127 ( .IN1(\R[0][0] ), .IN3(\R[2][0] ), .IN2(\R[1][0] ), .IN4(
        \R[3][0] ), .S0(N136), .S1(n7026), .Q(n6952) );
  MUX21X1 U6128 ( .IN1(n6952), .IN2(n6951), .S(N315), .Q(N594) );
  MUX41X1 U6129 ( .IN1(\R[4][1] ), .IN3(\R[6][1] ), .IN2(\R[5][1] ), .IN4(
        \R[7][1] ), .S0(N136), .S1(n7025), .Q(n6953) );
  MUX41X1 U6130 ( .IN1(\R[0][1] ), .IN3(\R[2][1] ), .IN2(\R[1][1] ), .IN4(
        \R[3][1] ), .S0(N136), .S1(n7025), .Q(n6954) );
  MUX21X1 U6131 ( .IN1(n6954), .IN2(n6953), .S(N315), .Q(N593) );
  MUX41X1 U6132 ( .IN1(\R[4][2] ), .IN3(\R[6][2] ), .IN2(\R[5][2] ), .IN4(
        \R[7][2] ), .S0(N136), .S1(n7018), .Q(n6955) );
  MUX41X1 U6133 ( .IN1(\R[0][2] ), .IN3(\R[2][2] ), .IN2(\R[1][2] ), .IN4(
        \R[3][2] ), .S0(N136), .S1(n7024), .Q(n6956) );
  MUX21X1 U6134 ( .IN1(n6956), .IN2(n6955), .S(N315), .Q(N592) );
  MUX41X1 U6135 ( .IN1(\R[4][3] ), .IN3(\R[6][3] ), .IN2(\R[5][3] ), .IN4(
        \R[7][3] ), .S0(N136), .S1(n7020), .Q(n6957) );
  MUX41X1 U6136 ( .IN1(\R[0][3] ), .IN3(\R[2][3] ), .IN2(\R[1][3] ), .IN4(
        \R[3][3] ), .S0(N136), .S1(n7023), .Q(n6958) );
  MUX21X1 U6137 ( .IN1(n6958), .IN2(n6957), .S(N315), .Q(N591) );
  MUX41X1 U6138 ( .IN1(\R[4][4] ), .IN3(\R[6][4] ), .IN2(\R[5][4] ), .IN4(
        \R[7][4] ), .S0(N136), .S1(n7020), .Q(n6959) );
  MUX41X1 U6139 ( .IN1(\R[0][4] ), .IN3(\R[2][4] ), .IN2(\R[1][4] ), .IN4(
        \R[3][4] ), .S0(N136), .S1(n7022), .Q(n6960) );
  MUX21X1 U6140 ( .IN1(n6960), .IN2(n6959), .S(N315), .Q(N590) );
  MUX41X1 U6141 ( .IN1(\R[4][5] ), .IN3(\R[6][5] ), .IN2(\R[5][5] ), .IN4(
        \R[7][5] ), .S0(N136), .S1(n7016), .Q(n6961) );
  MUX41X1 U6142 ( .IN1(\R[0][5] ), .IN3(\R[2][5] ), .IN2(\R[1][5] ), .IN4(
        \R[3][5] ), .S0(N136), .S1(n7021), .Q(n6962) );
  MUX21X1 U6143 ( .IN1(n6962), .IN2(n6961), .S(N315), .Q(N589) );
  MUX41X1 U6144 ( .IN1(\R[4][6] ), .IN3(\R[6][6] ), .IN2(\R[5][6] ), .IN4(
        \R[7][6] ), .S0(N136), .S1(n7018), .Q(n6963) );
  MUX41X1 U6145 ( .IN1(\R[0][6] ), .IN3(\R[2][6] ), .IN2(\R[1][6] ), .IN4(
        \R[3][6] ), .S0(N136), .S1(n7020), .Q(n6964) );
  MUX21X1 U6146 ( .IN1(n6964), .IN2(n6963), .S(N315), .Q(N588) );
  MUX41X1 U6147 ( .IN1(\R[4][7] ), .IN3(\R[6][7] ), .IN2(\R[5][7] ), .IN4(
        \R[7][7] ), .S0(N136), .S1(n7016), .Q(n6965) );
  MUX41X1 U6148 ( .IN1(\R[0][7] ), .IN3(\R[2][7] ), .IN2(\R[1][7] ), .IN4(
        \R[3][7] ), .S0(N136), .S1(n7019), .Q(n6966) );
  MUX21X1 U6149 ( .IN1(n6966), .IN2(n6965), .S(N315), .Q(N587) );
  MUX41X1 U6150 ( .IN1(\R[4][8] ), .IN3(\R[6][8] ), .IN2(\R[5][8] ), .IN4(
        \R[7][8] ), .S0(N136), .S1(n7021), .Q(n6967) );
  MUX41X1 U6151 ( .IN1(\R[0][8] ), .IN3(\R[2][8] ), .IN2(\R[1][8] ), .IN4(
        \R[3][8] ), .S0(N136), .S1(n7018), .Q(n6968) );
  MUX21X1 U6152 ( .IN1(n6968), .IN2(n6967), .S(N315), .Q(N586) );
  MUX41X1 U6153 ( .IN1(\R[4][9] ), .IN3(\R[6][9] ), .IN2(\R[5][9] ), .IN4(
        \R[7][9] ), .S0(N136), .S1(n7025), .Q(n6969) );
  MUX41X1 U6154 ( .IN1(\R[0][9] ), .IN3(\R[2][9] ), .IN2(\R[1][9] ), .IN4(
        \R[3][9] ), .S0(N136), .S1(n7017), .Q(n6970) );
  MUX21X1 U6155 ( .IN1(n6970), .IN2(n6969), .S(N315), .Q(N585) );
  MUX41X1 U6156 ( .IN1(\R[4][10] ), .IN3(\R[6][10] ), .IN2(\R[5][10] ), .IN4(
        \R[7][10] ), .S0(N136), .S1(n7018), .Q(n6971) );
  MUX41X1 U6157 ( .IN1(\R[0][10] ), .IN3(\R[2][10] ), .IN2(\R[1][10] ), .IN4(
        \R[3][10] ), .S0(N136), .S1(n7023), .Q(n6972) );
  MUX21X1 U6158 ( .IN1(n6972), .IN2(n6971), .S(N315), .Q(N584) );
  MUX41X1 U6159 ( .IN1(\R[4][11] ), .IN3(\R[6][11] ), .IN2(\R[5][11] ), .IN4(
        \R[7][11] ), .S0(N136), .S1(n7020), .Q(n6973) );
  MUX41X1 U6160 ( .IN1(\R[0][11] ), .IN3(\R[2][11] ), .IN2(\R[1][11] ), .IN4(
        \R[3][11] ), .S0(N136), .S1(n7020), .Q(n6974) );
  MUX21X1 U6161 ( .IN1(n6974), .IN2(n6973), .S(N315), .Q(N583) );
  MUX41X1 U6162 ( .IN1(\R[4][12] ), .IN3(\R[6][12] ), .IN2(\R[5][12] ), .IN4(
        \R[7][12] ), .S0(N136), .S1(n7017), .Q(n6975) );
  MUX41X1 U6163 ( .IN1(\R[0][12] ), .IN3(\R[2][12] ), .IN2(\R[1][12] ), .IN4(
        \R[3][12] ), .S0(N136), .S1(n7022), .Q(n6976) );
  MUX21X1 U6164 ( .IN1(n6976), .IN2(n6975), .S(N315), .Q(N582) );
  MUX41X1 U6165 ( .IN1(\R[4][13] ), .IN3(\R[6][13] ), .IN2(\R[5][13] ), .IN4(
        \R[7][13] ), .S0(N136), .S1(n7019), .Q(n6977) );
  MUX41X1 U6166 ( .IN1(\R[0][13] ), .IN3(\R[2][13] ), .IN2(\R[1][13] ), .IN4(
        \R[3][13] ), .S0(N136), .S1(n7024), .Q(n6978) );
  MUX21X1 U6167 ( .IN1(n6978), .IN2(n6977), .S(N315), .Q(N581) );
  MUX41X1 U6168 ( .IN1(\R[4][14] ), .IN3(\R[6][14] ), .IN2(\R[5][14] ), .IN4(
        \R[7][14] ), .S0(N136), .S1(n7022), .Q(n6979) );
  MUX41X1 U6169 ( .IN1(\R[0][14] ), .IN3(\R[2][14] ), .IN2(\R[1][14] ), .IN4(
        \R[3][14] ), .S0(N136), .S1(n7017), .Q(n6980) );
  MUX21X1 U6170 ( .IN1(n6980), .IN2(n6979), .S(N315), .Q(N580) );
  MUX41X1 U6171 ( .IN1(\R[4][15] ), .IN3(\R[6][15] ), .IN2(\R[5][15] ), .IN4(
        \R[7][15] ), .S0(N136), .S1(n7020), .Q(n6981) );
  MUX41X1 U6172 ( .IN1(\R[0][15] ), .IN3(\R[2][15] ), .IN2(\R[1][15] ), .IN4(
        \R[3][15] ), .S0(N136), .S1(n7016), .Q(n6982) );
  MUX21X1 U6173 ( .IN1(n6982), .IN2(n6981), .S(N315), .Q(N579) );
  MUX41X1 U6174 ( .IN1(\R[4][16] ), .IN3(\R[6][16] ), .IN2(\R[5][16] ), .IN4(
        \R[7][16] ), .S0(N136), .S1(n7015), .Q(n6983) );
  MUX41X1 U6175 ( .IN1(\R[0][16] ), .IN3(\R[2][16] ), .IN2(\R[1][16] ), .IN4(
        \R[3][16] ), .S0(N136), .S1(n7025), .Q(n6984) );
  MUX21X1 U6176 ( .IN1(n6984), .IN2(n6983), .S(N315), .Q(N578) );
  MUX41X1 U6177 ( .IN1(\R[4][17] ), .IN3(\R[6][17] ), .IN2(\R[5][17] ), .IN4(
        \R[7][17] ), .S0(N136), .S1(n7023), .Q(n6985) );
  MUX41X1 U6178 ( .IN1(\R[0][17] ), .IN3(\R[2][17] ), .IN2(\R[1][17] ), .IN4(
        \R[3][17] ), .S0(N136), .S1(n7015), .Q(n6986) );
  MUX21X1 U6179 ( .IN1(n6986), .IN2(n6985), .S(N315), .Q(N577) );
  MUX41X1 U6180 ( .IN1(\R[4][18] ), .IN3(\R[6][18] ), .IN2(\R[5][18] ), .IN4(
        \R[7][18] ), .S0(N136), .S1(n7022), .Q(n6987) );
  MUX41X1 U6181 ( .IN1(\R[0][18] ), .IN3(\R[2][18] ), .IN2(\R[1][18] ), .IN4(
        \R[3][18] ), .S0(N136), .S1(n7016), .Q(n6988) );
  MUX21X1 U6182 ( .IN1(n6988), .IN2(n6987), .S(N315), .Q(N576) );
  MUX41X1 U6183 ( .IN1(\R[4][19] ), .IN3(\R[6][19] ), .IN2(\R[5][19] ), .IN4(
        \R[7][19] ), .S0(N136), .S1(n7026), .Q(n6989) );
  MUX41X1 U6184 ( .IN1(\R[0][19] ), .IN3(\R[2][19] ), .IN2(\R[1][19] ), .IN4(
        \R[3][19] ), .S0(N136), .S1(n7015), .Q(n6990) );
  MUX21X1 U6185 ( .IN1(n6990), .IN2(n6989), .S(N315), .Q(N575) );
  MUX41X1 U6186 ( .IN1(\R[4][20] ), .IN3(\R[6][20] ), .IN2(\R[5][20] ), .IN4(
        \R[7][20] ), .S0(N136), .S1(n5697), .Q(n6991) );
  MUX41X1 U6187 ( .IN1(\R[0][20] ), .IN3(\R[2][20] ), .IN2(\R[1][20] ), .IN4(
        \R[3][20] ), .S0(N136), .S1(n7017), .Q(n6992) );
  MUX21X1 U6188 ( .IN1(n6992), .IN2(n6991), .S(N315), .Q(N574) );
  MUX41X1 U6189 ( .IN1(\R[4][21] ), .IN3(\R[6][21] ), .IN2(\R[5][21] ), .IN4(
        \R[7][21] ), .S0(N136), .S1(n7019), .Q(n6993) );
  MUX41X1 U6190 ( .IN1(\R[0][21] ), .IN3(\R[2][21] ), .IN2(\R[1][21] ), .IN4(
        \R[3][21] ), .S0(N136), .S1(n7016), .Q(n6994) );
  MUX21X1 U6191 ( .IN1(n6994), .IN2(n6993), .S(N315), .Q(N573) );
  MUX41X1 U6192 ( .IN1(\R[4][22] ), .IN3(\R[6][22] ), .IN2(\R[5][22] ), .IN4(
        \R[7][22] ), .S0(N136), .S1(n7018), .Q(n6995) );
  MUX41X1 U6193 ( .IN1(\R[0][22] ), .IN3(\R[2][22] ), .IN2(\R[1][22] ), .IN4(
        \R[3][22] ), .S0(N136), .S1(n7015), .Q(n6996) );
  MUX21X1 U6194 ( .IN1(n6996), .IN2(n6995), .S(N315), .Q(N572) );
  MUX41X1 U6195 ( .IN1(\R[4][23] ), .IN3(\R[6][23] ), .IN2(\R[5][23] ), .IN4(
        \R[7][23] ), .S0(N136), .S1(n5697), .Q(n6997) );
  MUX41X1 U6196 ( .IN1(\R[0][23] ), .IN3(\R[2][23] ), .IN2(\R[1][23] ), .IN4(
        \R[3][23] ), .S0(N136), .S1(n7017), .Q(n6998) );
  MUX21X1 U6197 ( .IN1(n6998), .IN2(n6997), .S(N315), .Q(N571) );
  MUX41X1 U6198 ( .IN1(\R[4][24] ), .IN3(\R[6][24] ), .IN2(\R[5][24] ), .IN4(
        \R[7][24] ), .S0(N136), .S1(n7019), .Q(n6999) );
  MUX41X1 U6199 ( .IN1(\R[0][24] ), .IN3(\R[2][24] ), .IN2(\R[1][24] ), .IN4(
        \R[3][24] ), .S0(N136), .S1(n7019), .Q(n7000) );
  MUX21X1 U6200 ( .IN1(n7000), .IN2(n6999), .S(N315), .Q(N570) );
  MUX41X1 U6201 ( .IN1(\R[4][25] ), .IN3(\R[6][25] ), .IN2(\R[5][25] ), .IN4(
        \R[7][25] ), .S0(N136), .S1(n7015), .Q(n7001) );
  MUX41X1 U6202 ( .IN1(\R[0][25] ), .IN3(\R[2][25] ), .IN2(\R[1][25] ), .IN4(
        \R[3][25] ), .S0(N136), .S1(n7024), .Q(n7002) );
  MUX21X1 U6203 ( .IN1(n7002), .IN2(n7001), .S(N315), .Q(N569) );
  MUX41X1 U6204 ( .IN1(\R[4][26] ), .IN3(\R[6][26] ), .IN2(\R[5][26] ), .IN4(
        \R[7][26] ), .S0(N136), .S1(n7024), .Q(n7003) );
  MUX41X1 U6205 ( .IN1(\R[0][26] ), .IN3(\R[2][26] ), .IN2(\R[1][26] ), .IN4(
        \R[3][26] ), .S0(N136), .S1(n7025), .Q(n7004) );
  MUX21X1 U6206 ( .IN1(n7004), .IN2(n7003), .S(N315), .Q(N568) );
  MUX41X1 U6207 ( .IN1(\R[4][27] ), .IN3(\R[6][27] ), .IN2(\R[5][27] ), .IN4(
        \R[7][27] ), .S0(N136), .S1(n7015), .Q(n7005) );
  MUX41X1 U6208 ( .IN1(\R[0][27] ), .IN3(\R[2][27] ), .IN2(\R[1][27] ), .IN4(
        \R[3][27] ), .S0(N136), .S1(n7023), .Q(n7006) );
  MUX21X1 U6209 ( .IN1(n7006), .IN2(n7005), .S(N315), .Q(N567) );
  MUX41X1 U6210 ( .IN1(\R[4][28] ), .IN3(\R[6][28] ), .IN2(\R[5][28] ), .IN4(
        \R[7][28] ), .S0(N136), .S1(n7024), .Q(n7007) );
  MUX41X1 U6211 ( .IN1(\R[0][28] ), .IN3(\R[2][28] ), .IN2(\R[1][28] ), .IN4(
        \R[3][28] ), .S0(N136), .S1(n7022), .Q(n7008) );
  MUX21X1 U6212 ( .IN1(n7008), .IN2(n7007), .S(N315), .Q(N566) );
  MUX41X1 U6213 ( .IN1(\R[4][29] ), .IN3(\R[6][29] ), .IN2(\R[5][29] ), .IN4(
        \R[7][29] ), .S0(N136), .S1(n7026), .Q(n7009) );
  MUX41X1 U6214 ( .IN1(\R[0][29] ), .IN3(\R[2][29] ), .IN2(\R[1][29] ), .IN4(
        \R[3][29] ), .S0(N136), .S1(n7016), .Q(n7010) );
  MUX21X1 U6215 ( .IN1(n7010), .IN2(n7009), .S(N315), .Q(N565) );
  MUX41X1 U6216 ( .IN1(\R[4][30] ), .IN3(\R[6][30] ), .IN2(\R[5][30] ), .IN4(
        \R[7][30] ), .S0(N136), .S1(n7023), .Q(n7011) );
  MUX41X1 U6217 ( .IN1(\R[0][30] ), .IN3(\R[2][30] ), .IN2(\R[1][30] ), .IN4(
        \R[3][30] ), .S0(N136), .S1(n7021), .Q(n7012) );
  MUX21X1 U6218 ( .IN1(n7012), .IN2(n7011), .S(N315), .Q(N564) );
  MUX41X1 U6219 ( .IN1(\R[4][31] ), .IN3(\R[6][31] ), .IN2(\R[5][31] ), .IN4(
        \R[7][31] ), .S0(N136), .S1(n5697), .Q(n7013) );
  MUX41X1 U6220 ( .IN1(\R[0][31] ), .IN3(\R[2][31] ), .IN2(\R[1][31] ), .IN4(
        \R[3][31] ), .S0(N136), .S1(n7026), .Q(n7014) );
  MUX21X1 U6221 ( .IN1(n7014), .IN2(n7013), .S(N315), .Q(N563) );
  MUX41X1 U6222 ( .IN1(\R[4][0] ), .IN3(\R[6][0] ), .IN2(\R[5][0] ), .IN4(
        \R[7][0] ), .S0(n5715), .S1(n5719), .Q(n7027) );
  MUX41X1 U6223 ( .IN1(\R[0][0] ), .IN3(\R[2][0] ), .IN2(\R[1][0] ), .IN4(
        \R[3][0] ), .S0(n5716), .S1(n5720), .Q(n7028) );
  MUX21X1 U6224 ( .IN1(n7028), .IN2(n7027), .S(N318), .Q(N5193) );
  MUX41X1 U6225 ( .IN1(\R[4][1] ), .IN3(\R[6][1] ), .IN2(\R[5][1] ), .IN4(
        \R[7][1] ), .S0(n5717), .S1(n5721), .Q(n7029) );
  MUX41X1 U6226 ( .IN1(\R[0][1] ), .IN3(\R[2][1] ), .IN2(\R[1][1] ), .IN4(
        \R[3][1] ), .S0(n5718), .S1(n5722), .Q(n7030) );
  MUX21X1 U6227 ( .IN1(n7030), .IN2(n7029), .S(N318), .Q(N5192) );
  MUX41X1 U6228 ( .IN1(\R[4][2] ), .IN3(\R[6][2] ), .IN2(\R[5][2] ), .IN4(
        \R[7][2] ), .S0(n5715), .S1(n5719), .Q(n7031) );
  MUX41X1 U6229 ( .IN1(\R[0][2] ), .IN3(\R[2][2] ), .IN2(\R[1][2] ), .IN4(
        \R[3][2] ), .S0(n5716), .S1(n5720), .Q(n7032) );
  MUX21X1 U6230 ( .IN1(n7032), .IN2(n7031), .S(N318), .Q(N5191) );
  MUX41X1 U6231 ( .IN1(\R[4][3] ), .IN3(\R[6][3] ), .IN2(\R[5][3] ), .IN4(
        \R[7][3] ), .S0(n5717), .S1(n5721), .Q(n7033) );
  MUX41X1 U6232 ( .IN1(\R[0][3] ), .IN3(\R[2][3] ), .IN2(\R[1][3] ), .IN4(
        \R[3][3] ), .S0(n5718), .S1(n5722), .Q(n7034) );
  MUX21X1 U6233 ( .IN1(n7034), .IN2(n7033), .S(N318), .Q(N5190) );
  MUX41X1 U6234 ( .IN1(\R[4][4] ), .IN3(\R[6][4] ), .IN2(\R[5][4] ), .IN4(
        \R[7][4] ), .S0(n5715), .S1(n5719), .Q(n7035) );
  MUX41X1 U6235 ( .IN1(\R[0][4] ), .IN3(\R[2][4] ), .IN2(\R[1][4] ), .IN4(
        \R[3][4] ), .S0(n5716), .S1(n5720), .Q(n7036) );
  MUX21X1 U6236 ( .IN1(n7036), .IN2(n7035), .S(N318), .Q(N5189) );
  MUX41X1 U6237 ( .IN1(\R[4][5] ), .IN3(\R[6][5] ), .IN2(\R[5][5] ), .IN4(
        \R[7][5] ), .S0(n5717), .S1(n5721), .Q(n7037) );
  MUX41X1 U6238 ( .IN1(\R[0][5] ), .IN3(\R[2][5] ), .IN2(\R[1][5] ), .IN4(
        \R[3][5] ), .S0(n5718), .S1(n5722), .Q(n7038) );
  MUX21X1 U6239 ( .IN1(n7038), .IN2(n7037), .S(N318), .Q(N5188) );
  MUX41X1 U6240 ( .IN1(\R[4][6] ), .IN3(\R[6][6] ), .IN2(\R[5][6] ), .IN4(
        \R[7][6] ), .S0(n5715), .S1(n5719), .Q(n7039) );
  MUX41X1 U6241 ( .IN1(\R[0][6] ), .IN3(\R[2][6] ), .IN2(\R[1][6] ), .IN4(
        \R[3][6] ), .S0(n5716), .S1(n5720), .Q(n7040) );
  MUX21X1 U6242 ( .IN1(n7040), .IN2(n7039), .S(N318), .Q(N5187) );
  MUX41X1 U6243 ( .IN1(\R[4][7] ), .IN3(\R[6][7] ), .IN2(\R[5][7] ), .IN4(
        \R[7][7] ), .S0(n5717), .S1(n5721), .Q(n7041) );
  MUX41X1 U6244 ( .IN1(\R[0][7] ), .IN3(\R[2][7] ), .IN2(\R[1][7] ), .IN4(
        \R[3][7] ), .S0(n5718), .S1(n5722), .Q(n7042) );
  MUX21X1 U6245 ( .IN1(n7042), .IN2(n7041), .S(N318), .Q(N5186) );
  MUX41X1 U6246 ( .IN1(\R[4][8] ), .IN3(\R[6][8] ), .IN2(\R[5][8] ), .IN4(
        \R[7][8] ), .S0(n5715), .S1(n5719), .Q(n7043) );
  MUX41X1 U6247 ( .IN1(\R[0][8] ), .IN3(\R[2][8] ), .IN2(\R[1][8] ), .IN4(
        \R[3][8] ), .S0(n5716), .S1(n5720), .Q(n7044) );
  MUX21X1 U6248 ( .IN1(n7044), .IN2(n7043), .S(N318), .Q(N5185) );
  MUX41X1 U6249 ( .IN1(\R[4][9] ), .IN3(\R[6][9] ), .IN2(\R[5][9] ), .IN4(
        \R[7][9] ), .S0(n5717), .S1(n5721), .Q(n7045) );
  MUX41X1 U6250 ( .IN1(\R[0][9] ), .IN3(\R[2][9] ), .IN2(\R[1][9] ), .IN4(
        \R[3][9] ), .S0(n5718), .S1(n5722), .Q(n7046) );
  MUX21X1 U6251 ( .IN1(n7046), .IN2(n7045), .S(N318), .Q(N5184) );
  MUX41X1 U6252 ( .IN1(\R[4][10] ), .IN3(\R[6][10] ), .IN2(\R[5][10] ), .IN4(
        \R[7][10] ), .S0(n5715), .S1(n5719), .Q(n7047) );
  MUX41X1 U6253 ( .IN1(\R[0][10] ), .IN3(\R[2][10] ), .IN2(\R[1][10] ), .IN4(
        \R[3][10] ), .S0(n5716), .S1(n5720), .Q(n7048) );
  MUX21X1 U6254 ( .IN1(n7048), .IN2(n7047), .S(N318), .Q(N5183) );
  MUX41X1 U6255 ( .IN1(\R[4][11] ), .IN3(\R[6][11] ), .IN2(\R[5][11] ), .IN4(
        \R[7][11] ), .S0(n5717), .S1(n5721), .Q(n7049) );
  MUX41X1 U6256 ( .IN1(\R[0][11] ), .IN3(\R[2][11] ), .IN2(\R[1][11] ), .IN4(
        \R[3][11] ), .S0(n5718), .S1(n5722), .Q(n7050) );
  MUX21X1 U6257 ( .IN1(n7050), .IN2(n7049), .S(N318), .Q(N5182) );
  MUX41X1 U6258 ( .IN1(\R[4][12] ), .IN3(\R[6][12] ), .IN2(\R[5][12] ), .IN4(
        \R[7][12] ), .S0(n5715), .S1(n5719), .Q(n7051) );
  MUX41X1 U6259 ( .IN1(\R[0][12] ), .IN3(\R[2][12] ), .IN2(\R[1][12] ), .IN4(
        \R[3][12] ), .S0(n5716), .S1(n5720), .Q(n7052) );
  MUX21X1 U6260 ( .IN1(n7052), .IN2(n7051), .S(N318), .Q(N5181) );
  MUX41X1 U6261 ( .IN1(\R[4][13] ), .IN3(\R[6][13] ), .IN2(\R[5][13] ), .IN4(
        \R[7][13] ), .S0(n5717), .S1(n5721), .Q(n7053) );
  MUX41X1 U6262 ( .IN1(\R[0][13] ), .IN3(\R[2][13] ), .IN2(\R[1][13] ), .IN4(
        \R[3][13] ), .S0(n5718), .S1(n5722), .Q(n7054) );
  MUX21X1 U6263 ( .IN1(n7054), .IN2(n7053), .S(N318), .Q(N5180) );
  MUX41X1 U6264 ( .IN1(\R[4][14] ), .IN3(\R[6][14] ), .IN2(\R[5][14] ), .IN4(
        \R[7][14] ), .S0(n5715), .S1(n5719), .Q(n7055) );
  MUX41X1 U6265 ( .IN1(\R[0][14] ), .IN3(\R[2][14] ), .IN2(\R[1][14] ), .IN4(
        \R[3][14] ), .S0(n5716), .S1(n5720), .Q(n7056) );
  MUX21X1 U6266 ( .IN1(n7056), .IN2(n7055), .S(N318), .Q(N5179) );
  MUX41X1 U6267 ( .IN1(\R[4][15] ), .IN3(\R[6][15] ), .IN2(\R[5][15] ), .IN4(
        \R[7][15] ), .S0(n5717), .S1(n5721), .Q(n7057) );
  MUX41X1 U6268 ( .IN1(\R[0][15] ), .IN3(\R[2][15] ), .IN2(\R[1][15] ), .IN4(
        \R[3][15] ), .S0(n5718), .S1(n5722), .Q(n7058) );
  MUX21X1 U6269 ( .IN1(n7058), .IN2(n7057), .S(N318), .Q(N5178) );
  MUX41X1 U6270 ( .IN1(\R[4][16] ), .IN3(\R[6][16] ), .IN2(\R[5][16] ), .IN4(
        \R[7][16] ), .S0(n5715), .S1(n5719), .Q(n7059) );
  MUX41X1 U6271 ( .IN1(\R[0][16] ), .IN3(\R[2][16] ), .IN2(\R[1][16] ), .IN4(
        \R[3][16] ), .S0(n5716), .S1(n5720), .Q(n7060) );
  MUX21X1 U6272 ( .IN1(n7060), .IN2(n7059), .S(N318), .Q(N5177) );
  MUX41X1 U6273 ( .IN1(\R[4][17] ), .IN3(\R[6][17] ), .IN2(\R[5][17] ), .IN4(
        \R[7][17] ), .S0(n5717), .S1(n5721), .Q(n7061) );
  MUX41X1 U6274 ( .IN1(\R[0][17] ), .IN3(\R[2][17] ), .IN2(\R[1][17] ), .IN4(
        \R[3][17] ), .S0(n5718), .S1(n5722), .Q(n7062) );
  MUX21X1 U6275 ( .IN1(n7062), .IN2(n7061), .S(N318), .Q(N5176) );
  MUX41X1 U6276 ( .IN1(\R[4][18] ), .IN3(\R[6][18] ), .IN2(\R[5][18] ), .IN4(
        \R[7][18] ), .S0(n5715), .S1(n5719), .Q(n7063) );
  MUX41X1 U6277 ( .IN1(\R[0][18] ), .IN3(\R[2][18] ), .IN2(\R[1][18] ), .IN4(
        \R[3][18] ), .S0(n5716), .S1(n5720), .Q(n7064) );
  MUX21X1 U6278 ( .IN1(n7064), .IN2(n7063), .S(N318), .Q(N5175) );
  MUX41X1 U6279 ( .IN1(\R[4][19] ), .IN3(\R[6][19] ), .IN2(\R[5][19] ), .IN4(
        \R[7][19] ), .S0(n5717), .S1(n5721), .Q(n7065) );
  MUX41X1 U6280 ( .IN1(\R[0][19] ), .IN3(\R[2][19] ), .IN2(\R[1][19] ), .IN4(
        \R[3][19] ), .S0(n5718), .S1(n5722), .Q(n7066) );
  MUX21X1 U6281 ( .IN1(n7066), .IN2(n7065), .S(N318), .Q(N5174) );
  MUX41X1 U6282 ( .IN1(\R[4][20] ), .IN3(\R[6][20] ), .IN2(\R[5][20] ), .IN4(
        \R[7][20] ), .S0(n5715), .S1(n5719), .Q(n7067) );
  MUX41X1 U6283 ( .IN1(\R[0][20] ), .IN3(\R[2][20] ), .IN2(\R[1][20] ), .IN4(
        \R[3][20] ), .S0(n5716), .S1(n5720), .Q(n7068) );
  MUX21X1 U6284 ( .IN1(n7068), .IN2(n7067), .S(N318), .Q(N5173) );
  MUX41X1 U6285 ( .IN1(\R[4][21] ), .IN3(\R[6][21] ), .IN2(\R[5][21] ), .IN4(
        \R[7][21] ), .S0(n5717), .S1(n5721), .Q(n7069) );
  MUX41X1 U6286 ( .IN1(\R[0][21] ), .IN3(\R[2][21] ), .IN2(\R[1][21] ), .IN4(
        \R[3][21] ), .S0(n5718), .S1(n5722), .Q(n7070) );
  MUX21X1 U6287 ( .IN1(n7070), .IN2(n7069), .S(N318), .Q(N5172) );
  MUX41X1 U6288 ( .IN1(\R[4][22] ), .IN3(\R[6][22] ), .IN2(\R[5][22] ), .IN4(
        \R[7][22] ), .S0(n5715), .S1(n5719), .Q(n7071) );
  MUX41X1 U6289 ( .IN1(\R[0][22] ), .IN3(\R[2][22] ), .IN2(\R[1][22] ), .IN4(
        \R[3][22] ), .S0(n5716), .S1(n5720), .Q(n7072) );
  MUX21X1 U6290 ( .IN1(n7072), .IN2(n7071), .S(N318), .Q(N5171) );
  MUX41X1 U6291 ( .IN1(\R[4][23] ), .IN3(\R[6][23] ), .IN2(\R[5][23] ), .IN4(
        \R[7][23] ), .S0(n5717), .S1(n5721), .Q(n7073) );
  MUX41X1 U6292 ( .IN1(\R[0][23] ), .IN3(\R[2][23] ), .IN2(\R[1][23] ), .IN4(
        \R[3][23] ), .S0(n5718), .S1(n5722), .Q(n7074) );
  MUX21X1 U6293 ( .IN1(n7074), .IN2(n7073), .S(N318), .Q(N5170) );
  MUX41X1 U6294 ( .IN1(\R[4][24] ), .IN3(\R[6][24] ), .IN2(\R[5][24] ), .IN4(
        \R[7][24] ), .S0(n5715), .S1(n5719), .Q(n7075) );
  MUX41X1 U6295 ( .IN1(\R[0][24] ), .IN3(\R[2][24] ), .IN2(\R[1][24] ), .IN4(
        \R[3][24] ), .S0(n5716), .S1(n5720), .Q(n7076) );
  MUX21X1 U6296 ( .IN1(n7076), .IN2(n7075), .S(N318), .Q(N5169) );
  MUX41X1 U6297 ( .IN1(\R[4][25] ), .IN3(\R[6][25] ), .IN2(\R[5][25] ), .IN4(
        \R[7][25] ), .S0(n5717), .S1(n5721), .Q(n7077) );
  MUX41X1 U6298 ( .IN1(\R[0][25] ), .IN3(\R[2][25] ), .IN2(\R[1][25] ), .IN4(
        \R[3][25] ), .S0(n5718), .S1(n5722), .Q(n7078) );
  MUX21X1 U6299 ( .IN1(n7078), .IN2(n7077), .S(N318), .Q(N5168) );
  MUX41X1 U6300 ( .IN1(\R[4][26] ), .IN3(\R[6][26] ), .IN2(\R[5][26] ), .IN4(
        \R[7][26] ), .S0(n5715), .S1(n5719), .Q(n7079) );
  MUX41X1 U6301 ( .IN1(\R[0][26] ), .IN3(\R[2][26] ), .IN2(\R[1][26] ), .IN4(
        \R[3][26] ), .S0(n5716), .S1(n5720), .Q(n7080) );
  MUX21X1 U6302 ( .IN1(n7080), .IN2(n7079), .S(N318), .Q(N5167) );
  MUX41X1 U6303 ( .IN1(\R[4][27] ), .IN3(\R[6][27] ), .IN2(\R[5][27] ), .IN4(
        \R[7][27] ), .S0(n5717), .S1(n5721), .Q(n7081) );
  MUX41X1 U6304 ( .IN1(\R[0][27] ), .IN3(\R[2][27] ), .IN2(\R[1][27] ), .IN4(
        \R[3][27] ), .S0(n5718), .S1(n5722), .Q(n7082) );
  MUX21X1 U6305 ( .IN1(n7082), .IN2(n7081), .S(N318), .Q(N5166) );
  MUX41X1 U6306 ( .IN1(\R[4][28] ), .IN3(\R[6][28] ), .IN2(\R[5][28] ), .IN4(
        \R[7][28] ), .S0(n5715), .S1(n5719), .Q(n7083) );
  MUX41X1 U6307 ( .IN1(\R[0][28] ), .IN3(\R[2][28] ), .IN2(\R[1][28] ), .IN4(
        \R[3][28] ), .S0(n5716), .S1(n5720), .Q(n7084) );
  MUX21X1 U6308 ( .IN1(n7084), .IN2(n7083), .S(N318), .Q(N5165) );
  MUX41X1 U6309 ( .IN1(\R[4][29] ), .IN3(\R[6][29] ), .IN2(\R[5][29] ), .IN4(
        \R[7][29] ), .S0(n5717), .S1(n5721), .Q(n7085) );
  MUX41X1 U6310 ( .IN1(\R[0][29] ), .IN3(\R[2][29] ), .IN2(\R[1][29] ), .IN4(
        \R[3][29] ), .S0(n5718), .S1(n5722), .Q(n7086) );
  MUX21X1 U6311 ( .IN1(n7086), .IN2(n7085), .S(N318), .Q(N5164) );
  MUX41X1 U6312 ( .IN1(\R[4][30] ), .IN3(\R[6][30] ), .IN2(\R[5][30] ), .IN4(
        \R[7][30] ), .S0(n5715), .S1(n5719), .Q(n7087) );
  MUX41X1 U6313 ( .IN1(\R[0][30] ), .IN3(\R[2][30] ), .IN2(\R[1][30] ), .IN4(
        \R[3][30] ), .S0(n5716), .S1(n5720), .Q(n7088) );
  MUX21X1 U6314 ( .IN1(n7088), .IN2(n7087), .S(N318), .Q(N5163) );
  MUX41X1 U6315 ( .IN1(\R[4][31] ), .IN3(\R[6][31] ), .IN2(\R[5][31] ), .IN4(
        \R[7][31] ), .S0(n5717), .S1(n5721), .Q(n7089) );
  MUX41X1 U6316 ( .IN1(\R[0][31] ), .IN3(\R[2][31] ), .IN2(\R[1][31] ), .IN4(
        \R[3][31] ), .S0(n5718), .S1(n5722), .Q(n7090) );
  MUX21X1 U6317 ( .IN1(n7090), .IN2(n7089), .S(N318), .Q(N5162) );
  OR2X1 U6318 ( .IN1(n7091), .IN2(n7092), .Q(n4421) );
  MUX21X1 U6319 ( .IN1(n425), .IN2(n9170), .S(n7093), .Q(n7091) );
  MUX21X1 U6320 ( .IN1(n9169), .IN2(n7094), .S(n7095), .Q(n4420) );
  NOR2X0 U6321 ( .IN1(n7096), .IN2(n7097), .QN(n7095) );
  OA21X1 U6322 ( .IN1(n7098), .IN2(n7099), .IN3(n7100), .Q(n7096) );
  XOR2X1 U6323 ( .IN1(n7101), .IN2(n7102), .Q(n7094) );
  OR2X1 U6324 ( .IN1(n7103), .IN2(n7104), .Q(n4418) );
  MUX21X1 U6325 ( .IN1(n7105), .IN2(instruction[9]), .S(reset_n), .Q(n7104) );
  OR2X1 U6326 ( .IN1(n7103), .IN2(n7106), .Q(n4417) );
  MUX21X1 U6327 ( .IN1(n7107), .IN2(instruction[10]), .S(reset_n), .Q(n7106)
         );
  OR2X1 U6328 ( .IN1(n7103), .IN2(n7108), .Q(n4416) );
  MUX21X1 U6329 ( .IN1(n9186), .IN2(instruction[11]), .S(reset_n), .Q(n7108)
         );
  OR2X1 U6330 ( .IN1(n7103), .IN2(n7109), .Q(n4415) );
  MUX21X1 U6331 ( .IN1(n9187), .IN2(instruction[12]), .S(reset_n), .Q(n7109)
         );
  OR2X1 U6332 ( .IN1(n7103), .IN2(n7110), .Q(n4414) );
  MUX21X1 U6333 ( .IN1(n9188), .IN2(instruction[14]), .S(reset_n), .Q(n7110)
         );
  OR2X1 U6334 ( .IN1(n7103), .IN2(n7111), .Q(n4413) );
  MUX21X1 U6335 ( .IN1(n9185), .IN2(instruction[15]), .S(reset_n), .Q(n7111)
         );
  INVX0 U6336 ( .INP(n7112), .ZN(n7103) );
  AO22X1 U6337 ( .IN1(n9189), .IN2(n7113), .IN3(instruction[13]), .IN4(n7114), 
        .Q(n4412) );
  MUX21X1 U6338 ( .IN1(ID_imm_offset[9]), .IN2(n7105), .S(n7115), .Q(n4411) );
  MUX21X1 U6339 ( .IN1(n7116), .IN2(n7107), .S(n7115), .Q(n4410) );
  AO22X1 U6340 ( .IN1(n9168), .IN2(n7117), .IN3(n7118), .IN4(n7105), .Q(n4409)
         );
  AO21X1 U6341 ( .IN1(n7119), .IN2(n7120), .IN3(n9168), .Q(n7118) );
  NAND2X0 U6342 ( .IN1(n9186), .IN2(n7107), .QN(n7120) );
  AO22X1 U6343 ( .IN1(n9190), .IN2(n7121), .IN3(n7119), .IN4(n7122), .Q(n4408)
         );
  AO21X1 U6344 ( .IN1(n7107), .IN2(n5702), .IN3(n7123), .Q(n7122) );
  NAND2X0 U6345 ( .IN1(n7119), .IN2(n4422), .QN(n7121) );
  NAND2X0 U6346 ( .IN1(n7124), .IN2(n7125), .QN(n4407) );
  OR3X1 U6347 ( .IN1(n5702), .IN2(n7126), .IN3(n7117), .Q(n7125) );
  OAI21X1 U6348 ( .IN1(n7117), .IN2(n9186), .IN3(n9167), .QN(n7124) );
  AO22X1 U6349 ( .IN1(n7021), .IN2(n7113), .IN3(instruction[8]), .IN4(n7114), 
        .Q(n4406) );
  MUX21X1 U6350 ( .IN1(n9166), .IN2(n7017), .S(n7127), .Q(n4405) );
  AND2X1 U6351 ( .IN1(n7128), .IN2(n7119), .Q(n7127) );
  INVX0 U6352 ( .INP(n7117), .ZN(n7119) );
  MUX21X1 U6353 ( .IN1(ID_imm_offset[8]), .IN2(n7019), .S(n7115), .Q(n4404) );
  AO22X1 U6354 ( .IN1(n7129), .IN2(n7113), .IN3(instruction[7]), .IN4(n7114), 
        .Q(n4403) );
  AO21X1 U6355 ( .IN1(n7130), .IN2(n7129), .IN3(n7131), .Q(n4402) );
  NOR4X0 U6356 ( .IN1(n3696), .IN2(n7115), .IN3(n7132), .IN4(n7133), .QN(n7131) );
  OA21X1 U6357 ( .IN1(n7134), .IN2(n5692), .IN3(n7135), .Q(n7133) );
  MUX21X1 U6358 ( .IN1(n7136), .IN2(n7137), .S(n9187), .Q(n7135) );
  NAND2X0 U6359 ( .IN1(n7138), .IN2(n7139), .QN(n7137) );
  XOR2X1 U6360 ( .IN1(n5686), .IN2(n9185), .Q(n7139) );
  NAND3X0 U6361 ( .IN1(n7140), .IN2(n7141), .IN3(n7142), .QN(n7136) );
  INVX0 U6362 ( .INP(n7143), .ZN(n7134) );
  NAND2X0 U6363 ( .IN1(n7144), .IN2(n7138), .QN(n7130) );
  OA22X1 U6364 ( .IN1(n7145), .IN2(n7146), .IN3(n7140), .IN4(n7147), .Q(n7138)
         );
  AO22X1 U6365 ( .IN1(n6947), .IN2(n7113), .IN3(instruction[6]), .IN4(n7114), 
        .Q(n4401) );
  MUX21X1 U6366 ( .IN1(n6945), .IN2(n7148), .S(n7149), .Q(n4400) );
  AO221X1 U6367 ( .IN1(N594), .IN2(n7150), .IN3(N498), .IN4(n7151), .IN5(n7152), .Q(n4399) );
  AO22X1 U6368 ( .IN1(N530), .IN2(n7153), .IN3(n7154), .IN4(n7155), .Q(n7152)
         );
  AO221X1 U6369 ( .IN1(N593), .IN2(n7150), .IN3(N497), .IN4(n7151), .IN5(n7156), .Q(n4398) );
  AO22X1 U6370 ( .IN1(N529), .IN2(n7153), .IN3(n7154), .IN4(n7157), .Q(n7156)
         );
  AO221X1 U6371 ( .IN1(N592), .IN2(n7150), .IN3(N496), .IN4(n7151), .IN5(n7158), .Q(n4397) );
  AO22X1 U6372 ( .IN1(N528), .IN2(n7153), .IN3(n7154), .IN4(n7159), .Q(n7158)
         );
  AO221X1 U6373 ( .IN1(N591), .IN2(n7150), .IN3(N495), .IN4(n7151), .IN5(n7160), .Q(n4396) );
  AO22X1 U6374 ( .IN1(N527), .IN2(n7153), .IN3(n7154), .IN4(n7161), .Q(n7160)
         );
  AO221X1 U6375 ( .IN1(N590), .IN2(n7150), .IN3(N494), .IN4(n7151), .IN5(n7162), .Q(n4395) );
  AO22X1 U6376 ( .IN1(N526), .IN2(n7153), .IN3(n7154), .IN4(n7163), .Q(n7162)
         );
  AO221X1 U6377 ( .IN1(N589), .IN2(n7150), .IN3(N493), .IN4(n7151), .IN5(n7164), .Q(n4394) );
  AO22X1 U6378 ( .IN1(N525), .IN2(n7153), .IN3(n7154), .IN4(n7165), .Q(n7164)
         );
  AO221X1 U6379 ( .IN1(N588), .IN2(n7150), .IN3(N492), .IN4(n7151), .IN5(n7166), .Q(n4393) );
  AO22X1 U6380 ( .IN1(N524), .IN2(n7153), .IN3(n7154), .IN4(n7167), .Q(n7166)
         );
  AO221X1 U6381 ( .IN1(N587), .IN2(n7150), .IN3(N491), .IN4(n7151), .IN5(n7168), .Q(n4392) );
  AO22X1 U6382 ( .IN1(N523), .IN2(n7153), .IN3(n7154), .IN4(n7169), .Q(n7168)
         );
  AO221X1 U6383 ( .IN1(N586), .IN2(n7150), .IN3(N490), .IN4(n7151), .IN5(n7170), .Q(n4391) );
  AO22X1 U6384 ( .IN1(N522), .IN2(n7153), .IN3(n7154), .IN4(n7171), .Q(n7170)
         );
  AO221X1 U6385 ( .IN1(N585), .IN2(n7150), .IN3(N489), .IN4(n7151), .IN5(n7172), .Q(n4390) );
  AO22X1 U6386 ( .IN1(N521), .IN2(n7153), .IN3(n7154), .IN4(n7173), .Q(n7172)
         );
  AO221X1 U6387 ( .IN1(N584), .IN2(n7150), .IN3(N488), .IN4(n7151), .IN5(n7174), .Q(n4389) );
  AO22X1 U6388 ( .IN1(N520), .IN2(n7153), .IN3(n7154), .IN4(n7175), .Q(n7174)
         );
  AO221X1 U6389 ( .IN1(N583), .IN2(n7150), .IN3(N487), .IN4(n7151), .IN5(n7176), .Q(n4388) );
  AO22X1 U6390 ( .IN1(N519), .IN2(n7153), .IN3(n7154), .IN4(n7177), .Q(n7176)
         );
  AO221X1 U6391 ( .IN1(N582), .IN2(n7150), .IN3(N486), .IN4(n7151), .IN5(n7178), .Q(n4387) );
  AO22X1 U6392 ( .IN1(N518), .IN2(n7153), .IN3(n7154), .IN4(n7179), .Q(n7178)
         );
  AO221X1 U6393 ( .IN1(N581), .IN2(n7150), .IN3(N485), .IN4(n7151), .IN5(n7180), .Q(n4386) );
  AO22X1 U6394 ( .IN1(N517), .IN2(n7153), .IN3(n7154), .IN4(n7181), .Q(n7180)
         );
  AO221X1 U6395 ( .IN1(N580), .IN2(n7150), .IN3(N484), .IN4(n7151), .IN5(n7182), .Q(n4385) );
  AO22X1 U6396 ( .IN1(N516), .IN2(n7153), .IN3(n7154), .IN4(n7183), .Q(n7182)
         );
  AO221X1 U6397 ( .IN1(N579), .IN2(n7150), .IN3(N483), .IN4(n7151), .IN5(n7184), .Q(n4384) );
  AO22X1 U6398 ( .IN1(N515), .IN2(n7153), .IN3(n7154), .IN4(n7185), .Q(n7184)
         );
  AO221X1 U6399 ( .IN1(N578), .IN2(n7150), .IN3(N482), .IN4(n7151), .IN5(n7186), .Q(n4383) );
  AO22X1 U6400 ( .IN1(N514), .IN2(n7153), .IN3(n7154), .IN4(n7187), .Q(n7186)
         );
  AO221X1 U6401 ( .IN1(N577), .IN2(n7150), .IN3(N481), .IN4(n7151), .IN5(n7188), .Q(n4382) );
  AO22X1 U6402 ( .IN1(N513), .IN2(n7153), .IN3(n7154), .IN4(n7189), .Q(n7188)
         );
  AO221X1 U6403 ( .IN1(N576), .IN2(n7150), .IN3(N480), .IN4(n7151), .IN5(n7190), .Q(n4381) );
  AO22X1 U6404 ( .IN1(N512), .IN2(n7153), .IN3(n7154), .IN4(n7191), .Q(n7190)
         );
  AO221X1 U6405 ( .IN1(N575), .IN2(n7150), .IN3(N479), .IN4(n7151), .IN5(n7192), .Q(n4380) );
  AO22X1 U6406 ( .IN1(N511), .IN2(n7153), .IN3(n7154), .IN4(n7193), .Q(n7192)
         );
  AO221X1 U6407 ( .IN1(N574), .IN2(n7150), .IN3(N478), .IN4(n7151), .IN5(n7194), .Q(n4379) );
  AO22X1 U6408 ( .IN1(N510), .IN2(n7153), .IN3(n7154), .IN4(n7195), .Q(n7194)
         );
  AO221X1 U6409 ( .IN1(N573), .IN2(n7150), .IN3(N477), .IN4(n7151), .IN5(n7196), .Q(n4378) );
  AO22X1 U6410 ( .IN1(N509), .IN2(n7153), .IN3(n7154), .IN4(n7197), .Q(n7196)
         );
  AO221X1 U6411 ( .IN1(N572), .IN2(n7150), .IN3(N476), .IN4(n7151), .IN5(n7198), .Q(n4377) );
  AO22X1 U6412 ( .IN1(N508), .IN2(n7153), .IN3(n7154), .IN4(n7199), .Q(n7198)
         );
  AO221X1 U6413 ( .IN1(N571), .IN2(n7150), .IN3(N475), .IN4(n7151), .IN5(n7200), .Q(n4376) );
  AO22X1 U6414 ( .IN1(N507), .IN2(n7153), .IN3(n7154), .IN4(n7201), .Q(n7200)
         );
  AO221X1 U6415 ( .IN1(N570), .IN2(n7150), .IN3(N474), .IN4(n7151), .IN5(n7202), .Q(n4375) );
  AO22X1 U6416 ( .IN1(N506), .IN2(n7153), .IN3(n7154), .IN4(n7203), .Q(n7202)
         );
  AO221X1 U6417 ( .IN1(N569), .IN2(n7150), .IN3(N473), .IN4(n7151), .IN5(n7204), .Q(n4374) );
  AO22X1 U6418 ( .IN1(N505), .IN2(n7153), .IN3(n7154), .IN4(n7205), .Q(n7204)
         );
  AO221X1 U6419 ( .IN1(N568), .IN2(n7150), .IN3(N472), .IN4(n7151), .IN5(n7206), .Q(n4373) );
  AO22X1 U6420 ( .IN1(N504), .IN2(n7153), .IN3(n7154), .IN4(n7207), .Q(n7206)
         );
  AO221X1 U6421 ( .IN1(N567), .IN2(n7150), .IN3(N471), .IN4(n7151), .IN5(n7208), .Q(n4372) );
  AO22X1 U6422 ( .IN1(N503), .IN2(n7153), .IN3(n7154), .IN4(n7209), .Q(n7208)
         );
  AO221X1 U6423 ( .IN1(N566), .IN2(n7150), .IN3(N470), .IN4(n7151), .IN5(n7210), .Q(n4371) );
  AO22X1 U6424 ( .IN1(N502), .IN2(n7153), .IN3(n7154), .IN4(n7211), .Q(n7210)
         );
  AO221X1 U6425 ( .IN1(N565), .IN2(n7150), .IN3(N469), .IN4(n7151), .IN5(n7212), .Q(n4370) );
  AO22X1 U6426 ( .IN1(N501), .IN2(n7153), .IN3(n7154), .IN4(n7213), .Q(n7212)
         );
  AO221X1 U6427 ( .IN1(N564), .IN2(n7150), .IN3(N468), .IN4(n7151), .IN5(n7214), .Q(n4369) );
  AO22X1 U6428 ( .IN1(N500), .IN2(n7153), .IN3(n7154), .IN4(n7215), .Q(n7214)
         );
  AO221X1 U6429 ( .IN1(N563), .IN2(n7150), .IN3(N467), .IN4(n7151), .IN5(n7216), .Q(n4368) );
  AO22X1 U6430 ( .IN1(N499), .IN2(n7153), .IN3(n7154), .IN4(n7217), .Q(n7216)
         );
  INVX0 U6431 ( .INP(n7218), .ZN(n7153) );
  NOR2X0 U6432 ( .IN1(n7219), .IN2(n7154), .QN(n7151) );
  INVX0 U6433 ( .INP(n7220), .ZN(n7154) );
  OA21X1 U6434 ( .IN1(n7221), .IN2(n7222), .IN3(n7220), .Q(n7150) );
  NAND4X0 U6435 ( .IN1(n7223), .IN2(n7218), .IN3(n7224), .IN4(n7225), .QN(
        n7220) );
  AOI21X1 U6436 ( .IN1(n7226), .IN2(n7227), .IN3(n7228), .QN(n7225) );
  NAND3X0 U6437 ( .IN1(n5686), .IN2(n5689), .IN3(n9185), .QN(n7224) );
  AO222X1 U6438 ( .IN1(n7229), .IN2(N563), .IN3(N499), .IN4(n7230), .IN5(n7231), .IN6(n7232), .Q(n4367) );
  AO222X1 U6439 ( .IN1(n7229), .IN2(N564), .IN3(N500), .IN4(n7230), .IN5(n7231), .IN6(n7233), .Q(n4366) );
  AO222X1 U6440 ( .IN1(n7229), .IN2(N565), .IN3(N501), .IN4(n7230), .IN5(n7231), .IN6(n7234), .Q(n4365) );
  AO222X1 U6441 ( .IN1(n7229), .IN2(N566), .IN3(N502), .IN4(n7230), .IN5(n7231), .IN6(n7235), .Q(n4364) );
  AO222X1 U6442 ( .IN1(n7229), .IN2(N567), .IN3(N503), .IN4(n7230), .IN5(n7231), .IN6(n7236), .Q(n4363) );
  AO222X1 U6443 ( .IN1(n7229), .IN2(N568), .IN3(N504), .IN4(n7230), .IN5(n7231), .IN6(n7237), .Q(n4362) );
  AO222X1 U6444 ( .IN1(n7229), .IN2(N569), .IN3(N505), .IN4(n7230), .IN5(n7231), .IN6(n7238), .Q(n4361) );
  AO222X1 U6445 ( .IN1(n7229), .IN2(N570), .IN3(N506), .IN4(n7230), .IN5(n7231), .IN6(n7239), .Q(n4360) );
  AO222X1 U6446 ( .IN1(n7229), .IN2(N571), .IN3(N507), .IN4(n7230), .IN5(n7231), .IN6(n7240), .Q(n4359) );
  AO222X1 U6447 ( .IN1(n7229), .IN2(N572), .IN3(N508), .IN4(n7230), .IN5(n7231), .IN6(n7241), .Q(n4358) );
  AO222X1 U6448 ( .IN1(n7229), .IN2(N573), .IN3(N509), .IN4(n7230), .IN5(n7231), .IN6(n7242), .Q(n4357) );
  AO222X1 U6449 ( .IN1(n7229), .IN2(N574), .IN3(N510), .IN4(n7230), .IN5(n7231), .IN6(n7243), .Q(n4356) );
  AO222X1 U6450 ( .IN1(n7229), .IN2(N575), .IN3(N511), .IN4(n7230), .IN5(n7231), .IN6(n7244), .Q(n4355) );
  AO222X1 U6451 ( .IN1(n7229), .IN2(N576), .IN3(N512), .IN4(n7230), .IN5(n7231), .IN6(n7245), .Q(n4354) );
  AO222X1 U6452 ( .IN1(n7229), .IN2(N577), .IN3(N513), .IN4(n7230), .IN5(n7231), .IN6(n7246), .Q(n4353) );
  AO222X1 U6453 ( .IN1(n7229), .IN2(N578), .IN3(N514), .IN4(n7230), .IN5(n7231), .IN6(n7247), .Q(n4352) );
  AO222X1 U6454 ( .IN1(n7229), .IN2(N579), .IN3(N515), .IN4(n7230), .IN5(n7231), .IN6(n7248), .Q(n4351) );
  AO222X1 U6455 ( .IN1(n7229), .IN2(N580), .IN3(N516), .IN4(n7230), .IN5(n7231), .IN6(n7249), .Q(n4350) );
  AO222X1 U6456 ( .IN1(n7229), .IN2(N581), .IN3(N517), .IN4(n7230), .IN5(n7231), .IN6(n7250), .Q(n4349) );
  AO222X1 U6457 ( .IN1(n7229), .IN2(N582), .IN3(N518), .IN4(n7230), .IN5(n7231), .IN6(n7251), .Q(n4348) );
  AO222X1 U6458 ( .IN1(n7229), .IN2(N583), .IN3(N519), .IN4(n7230), .IN5(n7231), .IN6(n7252), .Q(n4347) );
  AO222X1 U6459 ( .IN1(n7229), .IN2(N584), .IN3(N520), .IN4(n7230), .IN5(n7231), .IN6(n7253), .Q(n4346) );
  AO222X1 U6460 ( .IN1(n7229), .IN2(N585), .IN3(N521), .IN4(n7230), .IN5(n7231), .IN6(n7254), .Q(n4345) );
  AO222X1 U6461 ( .IN1(n7229), .IN2(N586), .IN3(N522), .IN4(n7230), .IN5(n7231), .IN6(n7255), .Q(n4344) );
  AO222X1 U6462 ( .IN1(n7229), .IN2(N587), .IN3(N523), .IN4(n7230), .IN5(n7231), .IN6(n7256), .Q(n4343) );
  AO222X1 U6463 ( .IN1(n7229), .IN2(N588), .IN3(N524), .IN4(n7230), .IN5(n7231), .IN6(n7257), .Q(n4342) );
  AO222X1 U6464 ( .IN1(n7229), .IN2(N589), .IN3(N525), .IN4(n7230), .IN5(n7231), .IN6(n7258), .Q(n4341) );
  AO222X1 U6465 ( .IN1(n7229), .IN2(N590), .IN3(N526), .IN4(n7230), .IN5(n7231), .IN6(n7259), .Q(n4340) );
  AO222X1 U6466 ( .IN1(n7229), .IN2(N591), .IN3(N527), .IN4(n7230), .IN5(n7231), .IN6(n7260), .Q(n4339) );
  AO222X1 U6467 ( .IN1(n7229), .IN2(N592), .IN3(N528), .IN4(n7230), .IN5(n7231), .IN6(n7261), .Q(n4338) );
  AO222X1 U6468 ( .IN1(n7229), .IN2(N593), .IN3(N529), .IN4(n7230), .IN5(n7231), .IN6(n7262), .Q(n4337) );
  AO222X1 U6469 ( .IN1(n7229), .IN2(N594), .IN3(N530), .IN4(n7230), .IN5(n7231), .IN6(n7263), .Q(n4336) );
  AO222X1 U6470 ( .IN1(n7264), .IN2(n7265), .IN3(N562), .IN4(n7266), .IN5(N498), .IN6(n7267), .Q(n4335) );
  AO222X1 U6471 ( .IN1(n7264), .IN2(n7268), .IN3(N561), .IN4(n7266), .IN5(N497), .IN6(n7267), .Q(n4334) );
  AO222X1 U6472 ( .IN1(n7264), .IN2(n7269), .IN3(N560), .IN4(n7266), .IN5(N496), .IN6(n7267), .Q(n4333) );
  AO222X1 U6473 ( .IN1(n7264), .IN2(n7270), .IN3(N559), .IN4(n7266), .IN5(N495), .IN6(n7267), .Q(n4332) );
  AO222X1 U6474 ( .IN1(n7264), .IN2(n7271), .IN3(N558), .IN4(n7266), .IN5(N494), .IN6(n7267), .Q(n4331) );
  AO222X1 U6475 ( .IN1(n7264), .IN2(n7272), .IN3(N557), .IN4(n7266), .IN5(N493), .IN6(n7267), .Q(n4330) );
  AO222X1 U6476 ( .IN1(n7264), .IN2(n7273), .IN3(N556), .IN4(n7266), .IN5(N492), .IN6(n7267), .Q(n4329) );
  AO222X1 U6477 ( .IN1(n7264), .IN2(n7274), .IN3(N555), .IN4(n7266), .IN5(N491), .IN6(n7267), .Q(n4328) );
  AO222X1 U6478 ( .IN1(n7264), .IN2(n7275), .IN3(N554), .IN4(n7266), .IN5(N490), .IN6(n7267), .Q(n4327) );
  AO222X1 U6479 ( .IN1(n7264), .IN2(n7276), .IN3(N553), .IN4(n7266), .IN5(N489), .IN6(n7267), .Q(n4326) );
  AO222X1 U6480 ( .IN1(n7264), .IN2(n7277), .IN3(N552), .IN4(n7266), .IN5(N488), .IN6(n7267), .Q(n4325) );
  AO222X1 U6481 ( .IN1(n7264), .IN2(n7278), .IN3(N551), .IN4(n7266), .IN5(N487), .IN6(n7267), .Q(n4324) );
  AO222X1 U6482 ( .IN1(n7264), .IN2(n7279), .IN3(N550), .IN4(n7266), .IN5(N486), .IN6(n7267), .Q(n4323) );
  AO222X1 U6483 ( .IN1(n7264), .IN2(n7280), .IN3(N549), .IN4(n7266), .IN5(N485), .IN6(n7267), .Q(n4322) );
  AO222X1 U6484 ( .IN1(n7264), .IN2(n7281), .IN3(N548), .IN4(n7266), .IN5(N484), .IN6(n7267), .Q(n4321) );
  AO222X1 U6485 ( .IN1(n7264), .IN2(n7282), .IN3(N547), .IN4(n7266), .IN5(N483), .IN6(n7267), .Q(n4320) );
  AO222X1 U6486 ( .IN1(n7264), .IN2(n7283), .IN3(N546), .IN4(n7266), .IN5(N482), .IN6(n7267), .Q(n4319) );
  AO222X1 U6487 ( .IN1(n7264), .IN2(n7284), .IN3(N545), .IN4(n7266), .IN5(N481), .IN6(n7267), .Q(n4318) );
  AO222X1 U6488 ( .IN1(n7264), .IN2(n7285), .IN3(N544), .IN4(n7266), .IN5(N480), .IN6(n7267), .Q(n4317) );
  AO222X1 U6489 ( .IN1(n7264), .IN2(n7286), .IN3(N543), .IN4(n7266), .IN5(N479), .IN6(n7267), .Q(n4316) );
  AO222X1 U6490 ( .IN1(n7264), .IN2(n7287), .IN3(N542), .IN4(n7266), .IN5(N478), .IN6(n7267), .Q(n4315) );
  AO222X1 U6491 ( .IN1(n7264), .IN2(n7288), .IN3(N541), .IN4(n7266), .IN5(N477), .IN6(n7267), .Q(n4314) );
  AO222X1 U6492 ( .IN1(n7264), .IN2(n7289), .IN3(N540), .IN4(n7266), .IN5(N476), .IN6(n7267), .Q(n4313) );
  AO222X1 U6493 ( .IN1(n7264), .IN2(n7290), .IN3(N539), .IN4(n7266), .IN5(N475), .IN6(n7267), .Q(n4312) );
  AO222X1 U6494 ( .IN1(n7264), .IN2(n7291), .IN3(N538), .IN4(n7266), .IN5(N474), .IN6(n7267), .Q(n4311) );
  AO222X1 U6495 ( .IN1(n7264), .IN2(n7292), .IN3(N537), .IN4(n7266), .IN5(N473), .IN6(n7267), .Q(n4310) );
  AO222X1 U6496 ( .IN1(n7264), .IN2(n7293), .IN3(N536), .IN4(n7266), .IN5(N472), .IN6(n7267), .Q(n4309) );
  AO222X1 U6497 ( .IN1(n7264), .IN2(n7294), .IN3(N535), .IN4(n7266), .IN5(N471), .IN6(n7267), .Q(n4308) );
  AO222X1 U6498 ( .IN1(n7264), .IN2(n7295), .IN3(N534), .IN4(n7266), .IN5(N470), .IN6(n7267), .Q(n4307) );
  AO222X1 U6499 ( .IN1(n7264), .IN2(n7296), .IN3(N533), .IN4(n7266), .IN5(N469), .IN6(n7267), .Q(n4306) );
  AO222X1 U6500 ( .IN1(n7264), .IN2(n7297), .IN3(N532), .IN4(n7266), .IN5(N468), .IN6(n7267), .Q(n4305) );
  AO222X1 U6501 ( .IN1(n7264), .IN2(n7298), .IN3(N531), .IN4(n7266), .IN5(N467), .IN6(n7267), .Q(n4304) );
  AND2X1 U6502 ( .IN1(n7299), .IN2(n7228), .Q(n7266) );
  NAND2X0 U6503 ( .IN1(n7300), .IN2(n7301), .QN(n7228) );
  INVX0 U6504 ( .INP(n7299), .ZN(n7264) );
  NAND3X0 U6505 ( .IN1(n7302), .IN2(n7301), .IN3(n7303), .QN(n7299) );
  INVX0 U6506 ( .INP(n7267), .ZN(n7303) );
  NAND3X0 U6507 ( .IN1(n7218), .IN2(n7304), .IN3(n7305), .QN(n7267) );
  NAND2X0 U6508 ( .IN1(n7306), .IN2(n7307), .QN(n7305) );
  NAND2X0 U6509 ( .IN1(n7308), .IN2(n7309), .QN(n7218) );
  NAND3X0 U6510 ( .IN1(n7310), .IN2(n7311), .IN3(n7312), .QN(n7309) );
  NAND2X0 U6511 ( .IN1(n7306), .IN2(n4422), .QN(n7302) );
  AO22X1 U6512 ( .IN1(n7313), .IN2(n7113), .IN3(instruction[5]), .IN4(n7114), 
        .Q(n4303) );
  MUX21X1 U6513 ( .IN1(n7313), .IN2(n7314), .S(n7149), .Q(n4302) );
  AND2X1 U6514 ( .IN1(n7315), .IN2(n7144), .Q(n7149) );
  AND2X1 U6515 ( .IN1(n7316), .IN2(n7317), .Q(n7144) );
  INVX0 U6516 ( .INP(n9195), .ZN(n7313) );
  AO22X1 U6517 ( .IN1(n7318), .IN2(n7113), .IN3(instruction[4]), .IN4(n7114), 
        .Q(n4301) );
  MUX21X1 U6518 ( .IN1(n7319), .IN2(n7320), .S(n7321), .Q(n4300) );
  AO22X1 U6519 ( .IN1(n7322), .IN2(n7107), .IN3(n7323), .IN4(n7318), .Q(n7320)
         );
  INVX0 U6520 ( .INP(n9196), .ZN(n7318) );
  AO22X1 U6521 ( .IN1(n5699), .IN2(n7113), .IN3(instruction[3]), .IN4(n7114), 
        .Q(n4299) );
  MUX21X1 U6522 ( .IN1(n7324), .IN2(n7325), .S(n7321), .Q(n4298) );
  AO22X1 U6523 ( .IN1(n7322), .IN2(n7105), .IN3(n7323), .IN4(n5699), .Q(n7325)
         );
  AO22X1 U6524 ( .IN1(n7326), .IN2(n7113), .IN3(instruction[2]), .IN4(n7114), 
        .Q(n4297) );
  AO222X1 U6525 ( .IN1(n7327), .IN2(n7326), .IN3(n7328), .IN4(n7025), .IN5(
        n7329), .IN6(n7330), .Q(n4296) );
  AO222X1 U6526 ( .IN1(n7229), .IN2(n7107), .IN3(n7230), .IN4(n7326), .IN5(
        n9165), .IN6(n7231), .Q(n4295) );
  INVX0 U6527 ( .INP(n9192), .ZN(n7326) );
  AO22X1 U6528 ( .IN1(n7331), .IN2(n7113), .IN3(instruction[1]), .IN4(n7114), 
        .Q(n4294) );
  AO222X1 U6529 ( .IN1(n7327), .IN2(n7331), .IN3(n7328), .IN4(n7129), .IN5(
        n7329), .IN6(n7332), .Q(n4293) );
  AO222X1 U6530 ( .IN1(n7229), .IN2(n7105), .IN3(n7230), .IN4(n7331), .IN5(
        n9164), .IN6(n7231), .Q(n4292) );
  INVX0 U6531 ( .INP(n9193), .ZN(n7331) );
  AO22X1 U6532 ( .IN1(n7333), .IN2(n7113), .IN3(instruction[0]), .IN4(n7114), 
        .Q(n4291) );
  AO222X1 U6533 ( .IN1(n7327), .IN2(n7333), .IN3(n7328), .IN4(n6948), .IN5(
        n7329), .IN6(n7334), .Q(n4290) );
  NOR2X0 U6534 ( .IN1(n7329), .IN2(n7335), .QN(n7328) );
  INVX0 U6535 ( .INP(n7336), .ZN(n7329) );
  AND2X1 U6536 ( .IN1(n7323), .IN2(n7336), .Q(n7327) );
  AO21X1 U6537 ( .IN1(n7337), .IN2(n7107), .IN3(n7321), .Q(n7336) );
  NAND4X0 U6538 ( .IN1(n7338), .IN2(n7315), .IN3(n7316), .IN4(n7339), .QN(
        n7321) );
  NAND2X0 U6539 ( .IN1(n7340), .IN2(n7307), .QN(n7339) );
  NOR4X0 U6540 ( .IN1(n7341), .IN2(n7222), .IN3(n7132), .IN4(n7115), .QN(n7316) );
  NOR2X0 U6541 ( .IN1(n7342), .IN2(n7226), .QN(n7115) );
  OA21X1 U6542 ( .IN1(n7015), .IN2(n7343), .IN3(n7221), .Q(n7132) );
  INVX0 U6543 ( .INP(n7344), .ZN(n7341) );
  OA22X1 U6544 ( .IN1(n7145), .IN2(n7345), .IN3(n7140), .IN4(n7147), .Q(n7315)
         );
  INVX0 U6545 ( .INP(n7346), .ZN(n7338) );
  NAND4X0 U6546 ( .IN1(n7347), .IN2(n7348), .IN3(n7142), .IN4(n7140), .QN(
        n7323) );
  AO21X1 U6547 ( .IN1(n5692), .IN2(n5689), .IN3(n5705), .Q(n7347) );
  AO222X1 U6548 ( .IN1(n7229), .IN2(n5697), .IN3(n7230), .IN4(n7333), .IN5(
        n9163), .IN6(n7231), .Q(n4289) );
  INVX0 U6549 ( .INP(n7349), .ZN(n7231) );
  INVX0 U6550 ( .INP(n9194), .ZN(n7333) );
  NAND3X0 U6551 ( .IN1(n7301), .IN2(n7304), .IN3(n7335), .QN(n7230) );
  INVX0 U6552 ( .INP(n7322), .ZN(n7335) );
  NAND3X0 U6553 ( .IN1(n7350), .IN2(n7223), .IN3(n7351), .QN(n7322) );
  NAND2X0 U6554 ( .IN1(n7340), .IN2(n5689), .QN(n7351) );
  AND2X1 U6555 ( .IN1(n7352), .IN2(n7349), .Q(n7229) );
  NAND4X0 U6556 ( .IN1(n7219), .IN2(n7344), .IN3(n7353), .IN4(n7304), .QN(
        n7349) );
  NAND2X0 U6557 ( .IN1(n7308), .IN2(n7354), .QN(n7304) );
  NAND4X0 U6558 ( .IN1(n7355), .IN2(n7356), .IN3(n7357), .IN4(n7358), .QN(
        n7354) );
  OA21X1 U6559 ( .IN1(n7359), .IN2(n7360), .IN3(n7361), .Q(n7358) );
  AO21X1 U6560 ( .IN1(n7362), .IN2(n7360), .IN3(n7363), .Q(n7357) );
  NAND2X0 U6561 ( .IN1(n7222), .IN2(n7364), .QN(n7353) );
  AND3X1 U6562 ( .IN1(n7223), .IN2(n7365), .IN3(n7301), .Q(n7219) );
  NAND2X0 U6563 ( .IN1(n7308), .IN2(n7366), .QN(n7301) );
  NAND4X0 U6564 ( .IN1(n7367), .IN2(n7368), .IN3(n7369), .IN4(n7370), .QN(
        n7366) );
  NOR2X0 U6565 ( .IN1(n7371), .IN2(n7372), .QN(n7369) );
  INVX0 U6566 ( .INP(n7147), .ZN(n7371) );
  NAND4X0 U6567 ( .IN1(n7317), .IN2(n7348), .IN3(n7143), .IN4(n7140), .QN(
        n7352) );
  NAND2X0 U6568 ( .IN1(n7373), .IN2(n9187), .QN(n7317) );
  NAND2X0 U6569 ( .IN1(n7374), .IN2(n7112), .QN(n4288) );
  MUX21X1 U6570 ( .IN1(n5703), .IN2(n3720), .S(reset_n), .Q(n7374) );
  NAND2X0 U6571 ( .IN1(n7375), .IN2(n7112), .QN(n4287) );
  MUX21X1 U6572 ( .IN1(n5693), .IN2(n3716), .S(reset_n), .Q(n7375) );
  NAND2X0 U6573 ( .IN1(n7376), .IN2(n7112), .QN(n4286) );
  MUX21X1 U6574 ( .IN1(n5688), .IN2(n3723), .S(reset_n), .Q(n7376) );
  NAND2X0 U6575 ( .IN1(n7377), .IN2(n7112), .QN(n4285) );
  MUX21X1 U6576 ( .IN1(n5708), .IN2(\r1720/A[3] ), .S(reset_n), .Q(n7377) );
  NAND2X0 U6577 ( .IN1(n7378), .IN2(n7112), .QN(n4284) );
  MUX21X1 U6578 ( .IN1(n5710), .IN2(n3719), .S(reset_n), .Q(n7378) );
  NAND2X0 U6579 ( .IN1(n7379), .IN2(n7112), .QN(n4283) );
  NAND2X0 U6580 ( .IN1(n9191), .IN2(reset_n), .QN(n7112) );
  MUX21X1 U6581 ( .IN1(n5707), .IN2(n3721), .S(reset_n), .Q(n7379) );
  MUX21X1 U6582 ( .IN1(n9162), .IN2(n9163), .S(n7114), .Q(n4282) );
  MUX21X1 U6583 ( .IN1(n9161), .IN2(n9164), .S(n7114), .Q(n4281) );
  MUX21X1 U6584 ( .IN1(n9160), .IN2(n9165), .S(n7114), .Q(n4280) );
  AO222X1 U6585 ( .IN1(n7380), .IN2(n7263), .IN3(N5193), .IN4(n7381), .IN5(
        n9199), .IN6(n7382), .Q(n4279) );
  AO222X1 U6586 ( .IN1(n7380), .IN2(n7262), .IN3(N5192), .IN4(n7381), .IN5(
        n9200), .IN6(n7382), .Q(n4278) );
  AO222X1 U6587 ( .IN1(n7380), .IN2(n7261), .IN3(N5191), .IN4(n7381), .IN5(
        n9201), .IN6(n7382), .Q(n4277) );
  AO222X1 U6588 ( .IN1(n7380), .IN2(n7260), .IN3(N5190), .IN4(n7381), .IN5(
        n9202), .IN6(n7382), .Q(n4276) );
  AO222X1 U6589 ( .IN1(n7380), .IN2(n7259), .IN3(N5189), .IN4(n7381), .IN5(
        n9203), .IN6(n7382), .Q(n4275) );
  AO222X1 U6590 ( .IN1(n7380), .IN2(n7258), .IN3(N5188), .IN4(n7381), .IN5(
        n9204), .IN6(n7382), .Q(n4274) );
  AO222X1 U6591 ( .IN1(n7380), .IN2(n7257), .IN3(N5187), .IN4(n7381), .IN5(
        n9205), .IN6(n7382), .Q(n4273) );
  AO222X1 U6592 ( .IN1(n7380), .IN2(n7256), .IN3(N5186), .IN4(n7381), .IN5(
        n9206), .IN6(n7382), .Q(n4272) );
  AO222X1 U6593 ( .IN1(n7380), .IN2(n7255), .IN3(N5185), .IN4(n7381), .IN5(
        n9207), .IN6(n7382), .Q(n4271) );
  AO222X1 U6594 ( .IN1(n7380), .IN2(n7254), .IN3(N5184), .IN4(n7381), .IN5(
        n9208), .IN6(n7382), .Q(n4270) );
  AO222X1 U6595 ( .IN1(n7380), .IN2(n7253), .IN3(N5183), .IN4(n7381), .IN5(
        n9209), .IN6(n7382), .Q(n4269) );
  AO222X1 U6596 ( .IN1(n7380), .IN2(n7252), .IN3(N5182), .IN4(n7381), .IN5(
        n9210), .IN6(n7382), .Q(n4268) );
  AO222X1 U6597 ( .IN1(n7380), .IN2(n7251), .IN3(N5181), .IN4(n7381), .IN5(
        n9211), .IN6(n7382), .Q(n4267) );
  AO222X1 U6598 ( .IN1(n7380), .IN2(n7250), .IN3(N5180), .IN4(n7381), .IN5(
        n9212), .IN6(n7382), .Q(n4266) );
  AO222X1 U6599 ( .IN1(n7380), .IN2(n7249), .IN3(N5179), .IN4(n7381), .IN5(
        n9213), .IN6(n7382), .Q(n4265) );
  AO222X1 U6600 ( .IN1(n7380), .IN2(n7248), .IN3(N5178), .IN4(n7381), .IN5(
        n9214), .IN6(n7382), .Q(n4264) );
  AO222X1 U6601 ( .IN1(n7380), .IN2(n7247), .IN3(N5177), .IN4(n7381), .IN5(
        n9215), .IN6(n7382), .Q(n4263) );
  AO222X1 U6602 ( .IN1(n7380), .IN2(n7246), .IN3(N5176), .IN4(n7381), .IN5(
        n9216), .IN6(n7382), .Q(n4262) );
  AO222X1 U6603 ( .IN1(n7380), .IN2(n7245), .IN3(N5175), .IN4(n7381), .IN5(
        n9217), .IN6(n7382), .Q(n4261) );
  AO222X1 U6604 ( .IN1(n7380), .IN2(n7244), .IN3(N5174), .IN4(n7381), .IN5(
        n9218), .IN6(n7382), .Q(n4260) );
  AO222X1 U6605 ( .IN1(n7380), .IN2(n7243), .IN3(N5173), .IN4(n7381), .IN5(
        n9219), .IN6(n7382), .Q(n4259) );
  AO222X1 U6606 ( .IN1(n7380), .IN2(n7242), .IN3(N5172), .IN4(n7381), .IN5(
        n9220), .IN6(n7382), .Q(n4258) );
  AO222X1 U6607 ( .IN1(n7380), .IN2(n7241), .IN3(N5171), .IN4(n7381), .IN5(
        n9221), .IN6(n7382), .Q(n4257) );
  AO222X1 U6608 ( .IN1(n7380), .IN2(n7240), .IN3(N5170), .IN4(n7381), .IN5(
        n9222), .IN6(n7382), .Q(n4256) );
  AO222X1 U6609 ( .IN1(n7380), .IN2(n7239), .IN3(N5169), .IN4(n7381), .IN5(
        n9223), .IN6(n7382), .Q(n4255) );
  AO222X1 U6610 ( .IN1(n7380), .IN2(n7238), .IN3(N5168), .IN4(n7381), .IN5(
        n9224), .IN6(n7382), .Q(n4254) );
  AO222X1 U6611 ( .IN1(n7380), .IN2(n7237), .IN3(N5167), .IN4(n7381), .IN5(
        n9225), .IN6(n7382), .Q(n4253) );
  AO222X1 U6612 ( .IN1(n7380), .IN2(n7236), .IN3(N5166), .IN4(n7381), .IN5(
        n9226), .IN6(n7382), .Q(n4252) );
  AO222X1 U6613 ( .IN1(n7380), .IN2(n7235), .IN3(N5165), .IN4(n7381), .IN5(
        n9227), .IN6(n7382), .Q(n4251) );
  AO222X1 U6614 ( .IN1(n7380), .IN2(n7234), .IN3(N5164), .IN4(n7381), .IN5(
        n9228), .IN6(n7382), .Q(n4250) );
  AO222X1 U6615 ( .IN1(n7380), .IN2(n7233), .IN3(N5163), .IN4(n7381), .IN5(
        n9229), .IN6(n7382), .Q(n4249) );
  AO222X1 U6616 ( .IN1(n7380), .IN2(n7232), .IN3(N5162), .IN4(n7381), .IN5(
        n9230), .IN6(n7382), .Q(n4248) );
  AND2X1 U6617 ( .IN1(n7383), .IN2(n7384), .Q(n7381) );
  NOR2X0 U6618 ( .IN1(n7384), .IN2(n7382), .QN(n7380) );
  INVX0 U6619 ( .INP(n7383), .ZN(n7382) );
  NOR2X0 U6620 ( .IN1(n7113), .IN2(N6325), .QN(n7383) );
  INVX0 U6621 ( .INP(reset_n), .ZN(n7113) );
  MUX21X1 U6622 ( .IN1(n7385), .IN2(n9174), .S(n7386), .Q(n4247) );
  MUX21X1 U6623 ( .IN1(n7148), .IN2(n9159), .S(n7386), .Q(n4246) );
  MUX21X1 U6624 ( .IN1(n7314), .IN2(n9175), .S(n7386), .Q(n4245) );
  MUX21X1 U6625 ( .IN1(n7319), .IN2(n9158), .S(n7386), .Q(n4244) );
  MUX21X1 U6626 ( .IN1(n7324), .IN2(n9178), .S(n7386), .Q(n4243) );
  MUX21X1 U6627 ( .IN1(n7330), .IN2(n9177), .S(n7386), .Q(n4242) );
  MUX21X1 U6628 ( .IN1(n7332), .IN2(n9176), .S(n7386), .Q(n4241) );
  AO222X1 U6629 ( .IN1(N1831), .IN2(n7387), .IN3(n507), .IN4(n7388), .IN5(
        n7389), .IN6(SP[31]), .Q(n4240) );
  AO222X1 U6630 ( .IN1(N1800), .IN2(n7387), .IN3(n538), .IN4(n7388), .IN5(
        n7389), .IN6(n7390), .Q(n4239) );
  AO222X1 U6631 ( .IN1(N1801), .IN2(n7387), .IN3(n537), .IN4(n7388), .IN5(
        n7389), .IN6(n7391), .Q(n4238) );
  AO222X1 U6632 ( .IN1(N1802), .IN2(n7387), .IN3(n536), .IN4(n7388), .IN5(
        n7389), .IN6(SP[2]), .Q(n4237) );
  AO222X1 U6633 ( .IN1(N1803), .IN2(n7387), .IN3(n535), .IN4(n7388), .IN5(
        n7389), .IN6(SP[3]), .Q(n4236) );
  AO222X1 U6634 ( .IN1(N1804), .IN2(n7387), .IN3(n534), .IN4(n7388), .IN5(
        n7389), .IN6(SP[4]), .Q(n4235) );
  AO222X1 U6635 ( .IN1(N1805), .IN2(n7387), .IN3(n533), .IN4(n7388), .IN5(
        n7389), .IN6(SP[5]), .Q(n4234) );
  AO222X1 U6636 ( .IN1(N1806), .IN2(n7387), .IN3(n532), .IN4(n7388), .IN5(
        n7389), .IN6(SP[6]), .Q(n4233) );
  AO222X1 U6637 ( .IN1(N1807), .IN2(n7387), .IN3(n531), .IN4(n7388), .IN5(
        n7389), .IN6(SP[7]), .Q(n4232) );
  AO222X1 U6638 ( .IN1(N1808), .IN2(n7387), .IN3(n530), .IN4(n7388), .IN5(
        n7389), .IN6(SP[8]), .Q(n4231) );
  AO222X1 U6639 ( .IN1(N1809), .IN2(n7387), .IN3(n529), .IN4(n7388), .IN5(
        n7389), .IN6(SP[9]), .Q(n4230) );
  AO222X1 U6640 ( .IN1(N1810), .IN2(n7387), .IN3(n528), .IN4(n7388), .IN5(
        n7389), .IN6(SP[10]), .Q(n4229) );
  AO222X1 U6641 ( .IN1(N1811), .IN2(n7387), .IN3(n527), .IN4(n7388), .IN5(
        n7389), .IN6(SP[11]), .Q(n4228) );
  AO222X1 U6642 ( .IN1(N1812), .IN2(n7387), .IN3(n526), .IN4(n7388), .IN5(
        n7389), .IN6(SP[12]), .Q(n4227) );
  AO222X1 U6643 ( .IN1(N1813), .IN2(n7387), .IN3(n525), .IN4(n7388), .IN5(
        n7389), .IN6(SP[13]), .Q(n4226) );
  AO222X1 U6644 ( .IN1(N1814), .IN2(n7387), .IN3(n524), .IN4(n7388), .IN5(
        n7389), .IN6(SP[14]), .Q(n4225) );
  AO222X1 U6645 ( .IN1(N1815), .IN2(n7387), .IN3(n523), .IN4(n7388), .IN5(
        n7389), .IN6(SP[15]), .Q(n4224) );
  AO222X1 U6646 ( .IN1(N1816), .IN2(n7387), .IN3(n522), .IN4(n7388), .IN5(
        n7389), .IN6(SP[16]), .Q(n4223) );
  AO222X1 U6647 ( .IN1(N1817), .IN2(n7387), .IN3(n521), .IN4(n7388), .IN5(
        n7389), .IN6(SP[17]), .Q(n4222) );
  AO222X1 U6648 ( .IN1(N1818), .IN2(n7387), .IN3(n520), .IN4(n7388), .IN5(
        n7389), .IN6(SP[18]), .Q(n4221) );
  AO222X1 U6649 ( .IN1(N1819), .IN2(n7387), .IN3(n519), .IN4(n7388), .IN5(
        n7389), .IN6(SP[19]), .Q(n4220) );
  AO222X1 U6650 ( .IN1(N1820), .IN2(n7387), .IN3(n518), .IN4(n7388), .IN5(
        n7389), .IN6(SP[20]), .Q(n4219) );
  AO222X1 U6651 ( .IN1(N1821), .IN2(n7387), .IN3(n517), .IN4(n7388), .IN5(
        n7389), .IN6(SP[21]), .Q(n4218) );
  AO222X1 U6652 ( .IN1(N1822), .IN2(n7387), .IN3(n516), .IN4(n7388), .IN5(
        n7389), .IN6(SP[22]), .Q(n4217) );
  AO222X1 U6653 ( .IN1(N1823), .IN2(n7387), .IN3(n515), .IN4(n7388), .IN5(
        n7389), .IN6(SP[23]), .Q(n4216) );
  AO222X1 U6654 ( .IN1(N1824), .IN2(n7387), .IN3(n514), .IN4(n7388), .IN5(
        n7389), .IN6(SP[24]), .Q(n4215) );
  AO222X1 U6655 ( .IN1(N1825), .IN2(n7387), .IN3(n513), .IN4(n7388), .IN5(
        n7389), .IN6(SP[25]), .Q(n4214) );
  AO222X1 U6656 ( .IN1(N1826), .IN2(n7387), .IN3(n512), .IN4(n7388), .IN5(
        n7389), .IN6(SP[26]), .Q(n4213) );
  AO222X1 U6657 ( .IN1(N1827), .IN2(n7387), .IN3(n511), .IN4(n7388), .IN5(
        n7389), .IN6(SP[27]), .Q(n4212) );
  AO222X1 U6658 ( .IN1(N1828), .IN2(n7387), .IN3(n510), .IN4(n7388), .IN5(
        n7389), .IN6(SP[28]), .Q(n4211) );
  AO222X1 U6659 ( .IN1(N1829), .IN2(n7387), .IN3(n509), .IN4(n7388), .IN5(
        n7389), .IN6(SP[29]), .Q(n4210) );
  AO222X1 U6660 ( .IN1(N1830), .IN2(n7387), .IN3(n508), .IN4(n7388), .IN5(
        n7389), .IN6(SP[30]), .Q(n4209) );
  AND2X1 U6661 ( .IN1(n7392), .IN2(n7393), .Q(n7388) );
  NAND3X0 U6662 ( .IN1(n7394), .IN2(n7395), .IN3(n3720), .QN(n7392) );
  NOR2X0 U6663 ( .IN1(n5753), .IN2(n7389), .QN(n7387) );
  INVX0 U6664 ( .INP(n7393), .ZN(n7389) );
  NAND3X0 U6665 ( .IN1(n7396), .IN2(n7386), .IN3(n7397), .QN(n7393) );
  NAND2X0 U6666 ( .IN1(n7398), .IN2(n3723), .QN(n7397) );
  NAND4X0 U6667 ( .IN1(n7399), .IN2(n7400), .IN3(n7401), .IN4(n7114), .QN(
        n7396) );
  MUX21X1 U6668 ( .IN1(n9157), .IN2(n7402), .S(n7403), .Q(n4208) );
  NOR2X0 U6669 ( .IN1(n7404), .IN2(n7097), .QN(n7403) );
  MUX21X1 U6670 ( .IN1(n9156), .IN2(N5622), .S(n7405), .Q(n4207) );
  AO221X1 U6671 ( .IN1(n7406), .IN2(N5622), .IN3(n7407), .IN4(n7390), .IN5(
        n7408), .Q(n4206) );
  AO22X1 U6672 ( .IN1(n7409), .IN2(data_address[0]), .IN3(n7410), .IN4(n538), 
        .Q(n7408) );
  MUX21X1 U6673 ( .IN1(n9155), .IN2(N5623), .S(n7405), .Q(n4205) );
  AO221X1 U6674 ( .IN1(N5623), .IN2(n7406), .IN3(n7407), .IN4(n7391), .IN5(
        n7411), .Q(n4204) );
  AO22X1 U6675 ( .IN1(n7409), .IN2(data_address[1]), .IN3(n7410), .IN4(n537), 
        .Q(n7411) );
  MUX21X1 U6676 ( .IN1(n9154), .IN2(N5624), .S(n7405), .Q(n4203) );
  AO221X1 U6677 ( .IN1(N5624), .IN2(n7406), .IN3(n7407), .IN4(SP[2]), .IN5(
        n7412), .Q(n4202) );
  AO22X1 U6678 ( .IN1(n7409), .IN2(data_address[2]), .IN3(n7410), .IN4(n536), 
        .Q(n7412) );
  MUX21X1 U6679 ( .IN1(n9153), .IN2(N5625), .S(n7405), .Q(n4201) );
  AO221X1 U6680 ( .IN1(N5625), .IN2(n7406), .IN3(n7407), .IN4(SP[3]), .IN5(
        n7413), .Q(n4200) );
  AO22X1 U6681 ( .IN1(n7409), .IN2(data_address[3]), .IN3(n7410), .IN4(n535), 
        .Q(n7413) );
  MUX21X1 U6682 ( .IN1(n9152), .IN2(N5626), .S(n7405), .Q(n4199) );
  AO221X1 U6683 ( .IN1(N5626), .IN2(n7406), .IN3(n7407), .IN4(SP[4]), .IN5(
        n7414), .Q(n4198) );
  AO22X1 U6684 ( .IN1(n7409), .IN2(data_address[4]), .IN3(n7410), .IN4(n534), 
        .Q(n7414) );
  MUX21X1 U6685 ( .IN1(n9151), .IN2(N5627), .S(n7405), .Q(n4197) );
  AO221X1 U6686 ( .IN1(N5627), .IN2(n7406), .IN3(n7407), .IN4(SP[5]), .IN5(
        n7415), .Q(n4196) );
  AO22X1 U6687 ( .IN1(n7409), .IN2(data_address[5]), .IN3(n7410), .IN4(n533), 
        .Q(n7415) );
  MUX21X1 U6688 ( .IN1(n9150), .IN2(N5628), .S(n7405), .Q(n4195) );
  AO221X1 U6689 ( .IN1(N5628), .IN2(n7406), .IN3(n7407), .IN4(SP[6]), .IN5(
        n7416), .Q(n4194) );
  AO22X1 U6690 ( .IN1(n7409), .IN2(data_address[6]), .IN3(n7410), .IN4(n532), 
        .Q(n7416) );
  MUX21X1 U6691 ( .IN1(n9149), .IN2(N5629), .S(n7405), .Q(n4193) );
  AO221X1 U6692 ( .IN1(N5629), .IN2(n7406), .IN3(n7407), .IN4(SP[7]), .IN5(
        n7417), .Q(n4192) );
  AO22X1 U6693 ( .IN1(n7409), .IN2(data_address[7]), .IN3(n7410), .IN4(n531), 
        .Q(n7417) );
  MUX21X1 U6694 ( .IN1(n9148), .IN2(N5630), .S(n7405), .Q(n4191) );
  AO221X1 U6695 ( .IN1(N5630), .IN2(n7406), .IN3(n7407), .IN4(SP[8]), .IN5(
        n7418), .Q(n4190) );
  AO22X1 U6696 ( .IN1(n7409), .IN2(data_address[8]), .IN3(n7410), .IN4(n530), 
        .Q(n7418) );
  MUX21X1 U6697 ( .IN1(n9147), .IN2(N5631), .S(n7405), .Q(n4189) );
  AO221X1 U6698 ( .IN1(N5631), .IN2(n7406), .IN3(n7407), .IN4(SP[9]), .IN5(
        n7419), .Q(n4188) );
  AO22X1 U6699 ( .IN1(n7409), .IN2(data_address[9]), .IN3(n7410), .IN4(n529), 
        .Q(n7419) );
  MUX21X1 U6700 ( .IN1(n9146), .IN2(N5632), .S(n7405), .Q(n4187) );
  AO221X1 U6701 ( .IN1(N5632), .IN2(n7406), .IN3(n7407), .IN4(SP[10]), .IN5(
        n7420), .Q(n4186) );
  AO22X1 U6702 ( .IN1(n7409), .IN2(data_address[10]), .IN3(n7410), .IN4(n528), 
        .Q(n7420) );
  MUX21X1 U6703 ( .IN1(n9145), .IN2(N5633), .S(n7405), .Q(n4185) );
  AO221X1 U6704 ( .IN1(N5633), .IN2(n7406), .IN3(n7407), .IN4(SP[11]), .IN5(
        n7421), .Q(n4184) );
  AO22X1 U6705 ( .IN1(n7409), .IN2(data_address[11]), .IN3(n7410), .IN4(n527), 
        .Q(n7421) );
  MUX21X1 U6706 ( .IN1(n9144), .IN2(N5634), .S(n7405), .Q(n4183) );
  AO221X1 U6707 ( .IN1(N5634), .IN2(n7406), .IN3(n7407), .IN4(SP[12]), .IN5(
        n7422), .Q(n4182) );
  AO22X1 U6708 ( .IN1(n7409), .IN2(data_address[12]), .IN3(n7410), .IN4(n526), 
        .Q(n7422) );
  MUX21X1 U6709 ( .IN1(n9143), .IN2(N5635), .S(n7405), .Q(n4181) );
  AO221X1 U6710 ( .IN1(N5635), .IN2(n7406), .IN3(n7407), .IN4(SP[13]), .IN5(
        n7423), .Q(n4180) );
  AO22X1 U6711 ( .IN1(n7409), .IN2(data_address[13]), .IN3(n7410), .IN4(n525), 
        .Q(n7423) );
  MUX21X1 U6712 ( .IN1(n9142), .IN2(N5636), .S(n7405), .Q(n4179) );
  AO221X1 U6713 ( .IN1(N5636), .IN2(n7406), .IN3(n7407), .IN4(SP[14]), .IN5(
        n7424), .Q(n4178) );
  AO22X1 U6714 ( .IN1(n7409), .IN2(data_address[14]), .IN3(n7410), .IN4(n524), 
        .Q(n7424) );
  MUX21X1 U6715 ( .IN1(n9141), .IN2(N5637), .S(n7405), .Q(n4177) );
  AO221X1 U6716 ( .IN1(N5637), .IN2(n7406), .IN3(n7407), .IN4(SP[15]), .IN5(
        n7425), .Q(n4176) );
  AO22X1 U6717 ( .IN1(n7409), .IN2(data_address[15]), .IN3(n7410), .IN4(n523), 
        .Q(n7425) );
  MUX21X1 U6718 ( .IN1(n9140), .IN2(N5638), .S(n7405), .Q(n4175) );
  AO221X1 U6719 ( .IN1(N5638), .IN2(n7406), .IN3(n7407), .IN4(SP[16]), .IN5(
        n7426), .Q(n4174) );
  AO22X1 U6720 ( .IN1(n7409), .IN2(data_address[16]), .IN3(n7410), .IN4(n522), 
        .Q(n7426) );
  MUX21X1 U6721 ( .IN1(n9139), .IN2(N5639), .S(n7405), .Q(n4173) );
  AO221X1 U6722 ( .IN1(N5639), .IN2(n7406), .IN3(n7407), .IN4(SP[17]), .IN5(
        n7427), .Q(n4172) );
  AO22X1 U6723 ( .IN1(n7409), .IN2(data_address[17]), .IN3(n7410), .IN4(n521), 
        .Q(n7427) );
  MUX21X1 U6724 ( .IN1(n9138), .IN2(N5640), .S(n7405), .Q(n4171) );
  AO221X1 U6725 ( .IN1(N5640), .IN2(n7406), .IN3(n7407), .IN4(SP[18]), .IN5(
        n7428), .Q(n4170) );
  AO22X1 U6726 ( .IN1(n7409), .IN2(data_address[18]), .IN3(n7410), .IN4(n520), 
        .Q(n7428) );
  MUX21X1 U6727 ( .IN1(n9137), .IN2(N5641), .S(n7405), .Q(n4169) );
  AO221X1 U6728 ( .IN1(N5641), .IN2(n7406), .IN3(n7407), .IN4(SP[19]), .IN5(
        n7429), .Q(n4168) );
  AO22X1 U6729 ( .IN1(n7409), .IN2(data_address[19]), .IN3(n7410), .IN4(n519), 
        .Q(n7429) );
  MUX21X1 U6730 ( .IN1(n9136), .IN2(N5642), .S(n7405), .Q(n4167) );
  AO221X1 U6731 ( .IN1(N5642), .IN2(n7406), .IN3(n7407), .IN4(SP[20]), .IN5(
        n7430), .Q(n4166) );
  AO22X1 U6732 ( .IN1(n7409), .IN2(data_address[20]), .IN3(n7410), .IN4(n518), 
        .Q(n7430) );
  MUX21X1 U6733 ( .IN1(n9135), .IN2(N5643), .S(n7405), .Q(n4165) );
  AO221X1 U6734 ( .IN1(N5643), .IN2(n7406), .IN3(n7407), .IN4(SP[21]), .IN5(
        n7431), .Q(n4164) );
  AO22X1 U6735 ( .IN1(n7409), .IN2(data_address[21]), .IN3(n7410), .IN4(n517), 
        .Q(n7431) );
  MUX21X1 U6736 ( .IN1(n9134), .IN2(N5644), .S(n7405), .Q(n4163) );
  AO221X1 U6737 ( .IN1(N5644), .IN2(n7406), .IN3(n7407), .IN4(SP[22]), .IN5(
        n7432), .Q(n4162) );
  AO22X1 U6738 ( .IN1(n7409), .IN2(data_address[22]), .IN3(n7410), .IN4(n516), 
        .Q(n7432) );
  MUX21X1 U6739 ( .IN1(n9133), .IN2(N5645), .S(n7405), .Q(n4161) );
  AO221X1 U6740 ( .IN1(N5645), .IN2(n7406), .IN3(n7407), .IN4(SP[23]), .IN5(
        n7433), .Q(n4160) );
  AO22X1 U6741 ( .IN1(n7409), .IN2(data_address[23]), .IN3(n7410), .IN4(n515), 
        .Q(n7433) );
  MUX21X1 U6742 ( .IN1(n9132), .IN2(N5646), .S(n7405), .Q(n4159) );
  AO221X1 U6743 ( .IN1(N5646), .IN2(n7406), .IN3(n7407), .IN4(SP[24]), .IN5(
        n7434), .Q(n4158) );
  AO22X1 U6744 ( .IN1(n7409), .IN2(data_address[24]), .IN3(n7410), .IN4(n514), 
        .Q(n7434) );
  MUX21X1 U6745 ( .IN1(n9131), .IN2(N5647), .S(n7405), .Q(n4157) );
  AO221X1 U6746 ( .IN1(N5647), .IN2(n7406), .IN3(n7407), .IN4(SP[25]), .IN5(
        n7435), .Q(n4156) );
  AO22X1 U6747 ( .IN1(n7409), .IN2(data_address[25]), .IN3(n7410), .IN4(n513), 
        .Q(n7435) );
  MUX21X1 U6748 ( .IN1(n9130), .IN2(N5648), .S(n7405), .Q(n4155) );
  AO221X1 U6749 ( .IN1(N5648), .IN2(n7406), .IN3(n7407), .IN4(SP[26]), .IN5(
        n7436), .Q(n4154) );
  AO22X1 U6750 ( .IN1(n7409), .IN2(data_address[26]), .IN3(n7410), .IN4(n512), 
        .Q(n7436) );
  MUX21X1 U6751 ( .IN1(n9129), .IN2(N5649), .S(n7405), .Q(n4153) );
  AO221X1 U6752 ( .IN1(N5649), .IN2(n7406), .IN3(n7407), .IN4(SP[27]), .IN5(
        n7437), .Q(n4152) );
  AO22X1 U6753 ( .IN1(n7409), .IN2(data_address[27]), .IN3(n7410), .IN4(n511), 
        .Q(n7437) );
  MUX21X1 U6754 ( .IN1(n9128), .IN2(N5650), .S(n7405), .Q(n4151) );
  AO221X1 U6755 ( .IN1(N5650), .IN2(n7406), .IN3(n7407), .IN4(SP[28]), .IN5(
        n7438), .Q(n4150) );
  AO22X1 U6756 ( .IN1(n7409), .IN2(data_address[28]), .IN3(n7410), .IN4(n510), 
        .Q(n7438) );
  MUX21X1 U6757 ( .IN1(n9127), .IN2(N5651), .S(n7405), .Q(n4149) );
  AO221X1 U6758 ( .IN1(N5651), .IN2(n7406), .IN3(n7407), .IN4(SP[29]), .IN5(
        n7439), .Q(n4148) );
  AO22X1 U6759 ( .IN1(n7409), .IN2(data_address[29]), .IN3(n7410), .IN4(n509), 
        .Q(n7439) );
  MUX21X1 U6760 ( .IN1(n9126), .IN2(N5652), .S(n7405), .Q(n4147) );
  AO221X1 U6761 ( .IN1(N5652), .IN2(n7406), .IN3(n7407), .IN4(SP[30]), .IN5(
        n7440), .Q(n4146) );
  AO22X1 U6762 ( .IN1(n7409), .IN2(data_address[30]), .IN3(n7410), .IN4(n508), 
        .Q(n7440) );
  NOR3X0 U6763 ( .IN1(n7441), .IN2(n7409), .IN3(n7442), .QN(n7406) );
  MUX21X1 U6764 ( .IN1(n9125), .IN2(N5653), .S(n7405), .Q(n4145) );
  AO221X1 U6765 ( .IN1(n7407), .IN2(SP[31]), .IN3(n7410), .IN4(n507), .IN5(
        n7443), .Q(n4144) );
  MUX21X1 U6766 ( .IN1(n7444), .IN2(data_address[31]), .S(n7409), .Q(n7443) );
  NOR2X0 U6767 ( .IN1(n7445), .IN2(n7442), .QN(n7444) );
  AND3X1 U6768 ( .IN1(n7442), .IN2(n7446), .IN3(n3716), .Q(n7410) );
  AND3X1 U6769 ( .IN1(n7446), .IN2(n7447), .IN3(n7442), .Q(n7407) );
  INVX0 U6770 ( .INP(n7409), .ZN(n7446) );
  OA21X1 U6771 ( .IN1(n7442), .IN2(n7097), .IN3(n7386), .Q(n7409) );
  NAND4X0 U6772 ( .IN1(n7448), .IN2(n7449), .IN3(n7450), .IN4(n7114), .QN(
        n7386) );
  MUX21X1 U6773 ( .IN1(n7451), .IN2(n7452), .S(n3716), .Q(n7448) );
  MUX21X1 U6774 ( .IN1(n7453), .IN2(n9124), .S(n7454), .Q(n4143) );
  MUX21X1 U6775 ( .IN1(n4424), .IN2(n7101), .S(n7455), .Q(n7453) );
  MUX21X1 U6776 ( .IN1(n7456), .IN2(n9123), .S(n7454), .Q(n4142) );
  AOI21X1 U6777 ( .IN1(n7114), .IN2(n7455), .IN3(n7398), .QN(n7454) );
  NOR3X0 U6778 ( .IN1(n7457), .IN2(n7097), .IN3(n7458), .QN(n7398) );
  NAND2X0 U6779 ( .IN1(n7459), .IN2(n7460), .QN(n7456) );
  NAND4X0 U6780 ( .IN1(n7461), .IN2(n7462), .IN3(n7463), .IN4(n7464), .QN(
        n7460) );
  NOR4X0 U6781 ( .IN1(n7465), .IN2(n7466), .IN3(n7467), .IN4(n7468), .QN(n7464) );
  OR4X1 U6782 ( .IN1(n7455), .IN2(N1254), .IN3(N1255), .IN4(n4424), .Q(n7468)
         );
  NOR2X0 U6783 ( .IN1(n3662), .IN2(n4454), .QN(n4424) );
  NAND2X0 U6784 ( .IN1(n7469), .IN2(n7470), .QN(n7455) );
  MUX21X1 U6785 ( .IN1(n7471), .IN2(n7472), .S(n7451), .Q(n7469) );
  NAND2X0 U6786 ( .IN1(n7450), .IN2(n3716), .QN(n7472) );
  OR4X1 U6787 ( .IN1(n4425), .IN2(n4426), .IN3(n4427), .IN4(n4428), .Q(n7467)
         );
  NOR2X0 U6788 ( .IN1(n3666), .IN2(n4458), .QN(n4428) );
  NOR2X0 U6789 ( .IN1(n3665), .IN2(n4457), .QN(n4427) );
  NOR2X0 U6790 ( .IN1(n3664), .IN2(n4456), .QN(n4426) );
  NOR2X0 U6791 ( .IN1(n3663), .IN2(n4455), .QN(n4425) );
  OR4X1 U6792 ( .IN1(n4429), .IN2(n4430), .IN3(n4431), .IN4(n4432), .Q(n7466)
         );
  NOR2X0 U6793 ( .IN1(n3670), .IN2(n4462), .QN(n4432) );
  NOR2X0 U6794 ( .IN1(n3669), .IN2(n4461), .QN(n4431) );
  NOR2X0 U6795 ( .IN1(n3668), .IN2(n4460), .QN(n4430) );
  NOR2X0 U6796 ( .IN1(n3667), .IN2(n4459), .QN(n4429) );
  OR4X1 U6797 ( .IN1(n4433), .IN2(n4434), .IN3(n4435), .IN4(n4436), .Q(n7465)
         );
  NOR2X0 U6798 ( .IN1(n3674), .IN2(n4466), .QN(n4436) );
  NOR2X0 U6799 ( .IN1(n3673), .IN2(n4465), .QN(n4435) );
  NOR2X0 U6800 ( .IN1(n3672), .IN2(n4464), .QN(n4434) );
  NOR2X0 U6801 ( .IN1(n3671), .IN2(n4463), .QN(n4433) );
  NOR4X0 U6802 ( .IN1(n7473), .IN2(n7474), .IN3(n4450), .IN4(n4449), .QN(n7463) );
  NOR2X0 U6803 ( .IN1(n3687), .IN2(n4479), .QN(n4449) );
  NOR2X0 U6804 ( .IN1(n3688), .IN2(n4480), .QN(n4450) );
  OR3X1 U6805 ( .IN1(n4452), .IN2(n4453), .IN3(n4451), .Q(n7474) );
  NOR2X0 U6806 ( .IN1(n3689), .IN2(n4481), .QN(n4451) );
  NOR2X0 U6807 ( .IN1(n3691), .IN2(n4483), .QN(n4453) );
  NOR2X0 U6808 ( .IN1(n3690), .IN2(n4482), .QN(n4452) );
  OR4X1 U6809 ( .IN1(n4445), .IN2(n4446), .IN3(n4447), .IN4(n4448), .Q(n7473)
         );
  NOR2X0 U6810 ( .IN1(n3686), .IN2(n4478), .QN(n4448) );
  NOR2X0 U6811 ( .IN1(n3685), .IN2(n4477), .QN(n4447) );
  NOR2X0 U6812 ( .IN1(n3684), .IN2(n4476), .QN(n4446) );
  NOR2X0 U6813 ( .IN1(n3683), .IN2(n4475), .QN(n4445) );
  NOR4X0 U6814 ( .IN1(n4444), .IN2(n4443), .IN3(n4442), .IN4(n4441), .QN(n7462) );
  NOR2X0 U6815 ( .IN1(n3679), .IN2(n4471), .QN(n4441) );
  NOR2X0 U6816 ( .IN1(n3680), .IN2(n4472), .QN(n4442) );
  NOR2X0 U6817 ( .IN1(n3681), .IN2(n4473), .QN(n4443) );
  NOR2X0 U6818 ( .IN1(n3682), .IN2(n4474), .QN(n4444) );
  NOR4X0 U6819 ( .IN1(n4440), .IN2(n4439), .IN3(n4438), .IN4(n4437), .QN(n7461) );
  NOR2X0 U6820 ( .IN1(n3675), .IN2(n4467), .QN(n4437) );
  NOR2X0 U6821 ( .IN1(n3676), .IN2(n4468), .QN(n4438) );
  NOR2X0 U6822 ( .IN1(n3677), .IN2(n4469), .QN(n4439) );
  NOR2X0 U6823 ( .IN1(n3678), .IN2(n4470), .QN(n4440) );
  NAND3X0 U6824 ( .IN1(n7445), .IN2(n7475), .IN3(n7476), .QN(n7459) );
  MUX21X1 U6825 ( .IN1(n7477), .IN2(n7478), .S(n7441), .Q(n7476) );
  NOR4X0 U6826 ( .IN1(n7479), .IN2(n7480), .IN3(n7481), .IN4(n7482), .QN(n7478) );
  OR4X1 U6827 ( .IN1(n9149), .IN2(n9148), .IN3(n9147), .IN4(n9146), .Q(n7482)
         );
  OR4X1 U6828 ( .IN1(n9145), .IN2(n9144), .IN3(n9143), .IN4(n9142), .Q(n7481)
         );
  OR4X1 U6829 ( .IN1(n9155), .IN2(n9154), .IN3(n9156), .IN4(n7483), .Q(n7480)
         );
  OR4X1 U6830 ( .IN1(n9150), .IN2(n9151), .IN3(n9152), .IN4(n9153), .Q(n7483)
         );
  OR4X1 U6831 ( .IN1(n7484), .IN2(n7485), .IN3(n7486), .IN4(n7487), .Q(n7479)
         );
  OR4X1 U6832 ( .IN1(n9133), .IN2(n9132), .IN3(n9131), .IN4(n9130), .Q(n7487)
         );
  OR4X1 U6833 ( .IN1(n9129), .IN2(n9128), .IN3(n9127), .IN4(n9126), .Q(n7486)
         );
  OR4X1 U6834 ( .IN1(n9141), .IN2(n9140), .IN3(n9139), .IN4(n9138), .Q(n7485)
         );
  OR4X1 U6835 ( .IN1(n9137), .IN2(n9136), .IN3(n9135), .IN4(n9134), .Q(n7484)
         );
  NOR4X0 U6836 ( .IN1(n7488), .IN2(n7489), .IN3(n7490), .IN4(n7491), .QN(n7477) );
  OR4X1 U6837 ( .IN1(N5629), .IN2(N5630), .IN3(N5631), .IN4(N5632), .Q(n7491)
         );
  OR4X1 U6838 ( .IN1(N5633), .IN2(N5634), .IN3(N5635), .IN4(N5636), .Q(n7490)
         );
  OR4X1 U6839 ( .IN1(N5623), .IN2(N5624), .IN3(N5622), .IN4(n7492), .Q(n7489)
         );
  OR4X1 U6840 ( .IN1(N5628), .IN2(N5627), .IN3(N5626), .IN4(N5625), .Q(n7492)
         );
  OR4X1 U6841 ( .IN1(n7493), .IN2(n7494), .IN3(n7495), .IN4(n7496), .Q(n7488)
         );
  OR4X1 U6842 ( .IN1(N5645), .IN2(N5646), .IN3(N5647), .IN4(N5648), .Q(n7496)
         );
  OR4X1 U6843 ( .IN1(N5649), .IN2(N5650), .IN3(N5651), .IN4(N5652), .Q(n7495)
         );
  OR4X1 U6844 ( .IN1(N5637), .IN2(N5638), .IN3(N5639), .IN4(N5640), .Q(n7494)
         );
  OR4X1 U6845 ( .IN1(N5641), .IN2(N5642), .IN3(N5643), .IN4(N5644), .Q(n7493)
         );
  NAND4X0 U6846 ( .IN1(n7100), .IN2(n7497), .IN3(n7498), .IN4(n7499), .QN(
        n7475) );
  NOR2X0 U6847 ( .IN1(n7500), .IN2(n7501), .QN(n7498) );
  AND4X1 U6848 ( .IN1(n7502), .IN2(n7503), .IN3(n7504), .IN4(n7505), .Q(n7100)
         );
  OA22X1 U6849 ( .IN1(n7506), .IN2(n3723), .IN3(n7457), .IN4(n7507), .Q(n7505)
         );
  NAND2X0 U6850 ( .IN1(n7500), .IN2(n3716), .QN(n7507) );
  OA21X1 U6851 ( .IN1(n7457), .IN2(n7508), .IN3(n7509), .Q(n7506) );
  NAND3X0 U6852 ( .IN1(n3721), .IN2(n7510), .IN3(n7511), .QN(n7502) );
  AO21X1 U6853 ( .IN1(n3723), .IN2(n7512), .IN3(n7513), .Q(n7510) );
  INVX0 U6854 ( .INP(n7101), .ZN(n7445) );
  MUX21X1 U6855 ( .IN1(n9173), .IN2(n7514), .S(n7515), .Q(n4141) );
  NOR2X0 U6856 ( .IN1(n7516), .IN2(n7097), .QN(n7515) );
  AND3X1 U6857 ( .IN1(n7517), .IN2(n7518), .IN3(n7519), .Q(n7516) );
  OA221X1 U6858 ( .IN1(n7520), .IN2(n7521), .IN3(n7499), .IN4(n7522), .IN5(
        n7523), .Q(n7519) );
  NAND4X0 U6859 ( .IN1(n7524), .IN2(n7450), .IN3(n7525), .IN4(n7526), .QN(
        n7523) );
  NAND2X0 U6860 ( .IN1(n7527), .IN2(n7528), .QN(n7525) );
  NAND2X0 U6861 ( .IN1(n7401), .IN2(n7529), .QN(n7522) );
  OA22X1 U6862 ( .IN1(n7499), .IN2(n7497), .IN3(n7530), .IN4(n7531), .Q(n7520)
         );
  NAND2X0 U6863 ( .IN1(n7532), .IN2(n7513), .QN(n7518) );
  AO22X1 U6864 ( .IN1(n7102), .IN2(n7533), .IN3(n7101), .IN4(n7534), .Q(n7514)
         );
  AO22X1 U6865 ( .IN1(n7527), .IN2(n7524), .IN3(n7535), .IN4(n7536), .Q(n7534)
         );
  INVX0 U6866 ( .INP(n7537), .ZN(n7535) );
  NAND3X0 U6867 ( .IN1(n7538), .IN2(n7517), .IN3(n7539), .QN(n7533) );
  OA221X1 U6868 ( .IN1(n7527), .IN2(n7540), .IN3(n7536), .IN4(n7537), .IN5(
        n7503), .Q(n7539) );
  OR2X1 U6869 ( .IN1(n7099), .IN2(n3723), .Q(n7503) );
  NAND2X0 U6870 ( .IN1(n7511), .IN2(n7401), .QN(n7099) );
  NAND3X0 U6871 ( .IN1(\r1720/A[3] ), .IN2(n5753), .IN3(n7511), .QN(n7537) );
  AND3X1 U6872 ( .IN1(n7541), .IN2(n7504), .IN3(n7542), .Q(n7517) );
  AO21X1 U6873 ( .IN1(n7543), .IN2(n7544), .IN3(n3716), .Q(n7504) );
  NAND2X0 U6874 ( .IN1(n7450), .IN2(n7500), .QN(n7543) );
  NAND3X0 U6875 ( .IN1(n7545), .IN2(n7447), .IN3(n7400), .QN(n7541) );
  MUX21X1 U6876 ( .IN1(n7402), .IN2(n9157), .S(n7404), .Q(n7102) );
  AND4X1 U6877 ( .IN1(n7546), .IN2(n7547), .IN3(n7548), .IN4(n7549), .Q(n7404)
         );
  NAND2X0 U6878 ( .IN1(n7511), .IN2(n7550), .QN(n7548) );
  MUX21X1 U6879 ( .IN1(n7551), .IN2(n7552), .S(n3719), .Q(n7547) );
  AOI21X1 U6880 ( .IN1(n7530), .IN2(n7452), .IN3(n7512), .QN(n7552) );
  NAND2X0 U6881 ( .IN1(n7499), .IN2(n7530), .QN(n7551) );
  MUX21X1 U6882 ( .IN1(n7553), .IN2(n7554), .S(\r1720/A[3] ), .Q(n7546) );
  NAND2X0 U6883 ( .IN1(n7555), .IN2(n7457), .QN(n7554) );
  OA22X1 U6884 ( .IN1(n7450), .IN2(n7556), .IN3(n5696), .IN4(n7499), .Q(n7553)
         );
  NAND4X0 U6885 ( .IN1(n7557), .IN2(n7558), .IN3(n7559), .IN4(n7560), .QN(
        n7402) );
  NOR3X0 U6886 ( .IN1(n7561), .IN2(n7562), .IN3(n7563), .QN(n7560) );
  MUX21X1 U6887 ( .IN1(n7564), .IN2(n7565), .S(\r1720/A[3] ), .Q(n7563) );
  NAND4X0 U6888 ( .IN1(n7566), .IN2(n7567), .IN3(n7568), .IN4(n7569), .QN(
        n7565) );
  OA22X1 U6889 ( .IN1(n7570), .IN2(n7499), .IN3(n7571), .IN4(n7447), .Q(n7569)
         );
  AOI22X1 U6890 ( .IN1(n7572), .IN2(N1767), .IN3(N4879), .IN4(n7450), .QN(
        n7571) );
  NOR2X0 U6891 ( .IN1(n7457), .IN2(n7556), .QN(n7572) );
  OA22X1 U6892 ( .IN1(n7573), .IN2(n7574), .IN3(n7457), .IN4(n7575), .Q(n7570)
         );
  INVX0 U6893 ( .INP(N4710), .ZN(n7575) );
  NAND2X0 U6894 ( .IN1(n7576), .IN2(n3719), .QN(n7574) );
  NAND3X0 U6895 ( .IN1(n7450), .IN2(n5695), .IN3(N4611), .QN(n7568) );
  NAND3X0 U6896 ( .IN1(n7524), .IN2(n3721), .IN3(N4776), .QN(n7567) );
  NAND3X0 U6897 ( .IN1(n7577), .IN2(n3720), .IN3(n393), .QN(n7566) );
  NOR2X0 U6898 ( .IN1(n7578), .IN2(n7579), .QN(n7564) );
  AOI221X1 U6899 ( .IN1(n7580), .IN2(n7581), .IN3(n7582), .IN4(n7583), .IN5(
        n7584), .QN(n7578) );
  AO222X1 U6900 ( .IN1(n7585), .IN2(n7586), .IN3(n7587), .IN4(n7588), .IN5(
        n7589), .IN6(n7590), .Q(n7582) );
  AO222X1 U6901 ( .IN1(n7591), .IN2(n7592), .IN3(n7593), .IN4(n7594), .IN5(
        n7595), .IN6(n7596), .Q(n7587) );
  AO221X1 U6902 ( .IN1(n7597), .IN2(n7598), .IN3(n7599), .IN4(n7600), .IN5(
        n7601), .Q(n7593) );
  OAI22X1 U6903 ( .IN1(n7602), .IN2(n7603), .IN3(n7604), .IN4(n7605), .QN(
        n7601) );
  AOI22X1 U6904 ( .IN1(n7606), .IN2(n7607), .IN3(n7608), .IN4(n7609), .QN(
        n7604) );
  AOI222X1 U6905 ( .IN1(n7610), .IN2(n7611), .IN3(n7612), .IN4(n7613), .IN5(
        n7614), .IN6(n7615), .QN(n7602) );
  AO222X1 U6906 ( .IN1(n7616), .IN2(n7617), .IN3(n7618), .IN4(n7619), .IN5(
        n7620), .IN6(n7621), .Q(n7612) );
  AO222X1 U6907 ( .IN1(n7622), .IN2(n7623), .IN3(n7624), .IN4(n7625), .IN5(
        n7626), .IN6(n7627), .Q(n7618) );
  AO222X1 U6908 ( .IN1(n7628), .IN2(n7629), .IN3(n7630), .IN4(n7631), .IN5(
        n7632), .IN6(n7633), .Q(n7624) );
  AO222X1 U6909 ( .IN1(n7634), .IN2(n7635), .IN3(n7636), .IN4(n7637), .IN5(
        n7638), .IN6(n7639), .Q(n7630) );
  AO222X1 U6910 ( .IN1(n7640), .IN2(n7641), .IN3(n7642), .IN4(n7643), .IN5(
        n7644), .IN6(n7645), .Q(n7636) );
  AO222X1 U6911 ( .IN1(n7646), .IN2(n7647), .IN3(n7648), .IN4(n7649), .IN5(
        n7650), .IN6(n7651), .Q(n7642) );
  AO222X1 U6912 ( .IN1(n7652), .IN2(n7653), .IN3(n7654), .IN4(n7655), .IN5(
        n7656), .IN6(n7657), .Q(n7648) );
  AO221X1 U6913 ( .IN1(n7658), .IN2(n7659), .IN3(n7660), .IN4(n7661), .IN5(
        n7662), .Q(n7654) );
  OAI22X1 U6914 ( .IN1(n7663), .IN2(n7664), .IN3(n7665), .IN4(n7666), .QN(
        n7662) );
  AOI22X1 U6915 ( .IN1(n7667), .IN2(n7668), .IN3(n7669), .IN4(n7670), .QN(
        n7665) );
  AOI22X1 U6916 ( .IN1(n7262), .IN2(n7671), .IN3(n7263), .IN4(n7672), .QN(
        n7663) );
  MUX21X1 U6917 ( .IN1(n7673), .IN2(n7674), .S(n3720), .Q(n7562) );
  NOR2X0 U6918 ( .IN1(n7675), .IN2(n7458), .QN(n7674) );
  AND3X1 U6919 ( .IN1(n7676), .IN2(n7677), .IN3(n7678), .Q(n7675) );
  MUX21X1 U6920 ( .IN1(n7679), .IN2(n7680), .S(n7681), .Q(n7678) );
  AOI222X1 U6921 ( .IN1(n7682), .IN2(n7683), .IN3(n7684), .IN4(n7685), .IN5(
        n7599), .IN6(n7686), .QN(n7680) );
  AO22X1 U6922 ( .IN1(n7687), .IN2(n7688), .IN3(n7689), .IN4(n7690), .Q(n7685)
         );
  INVX0 U6923 ( .INP(n7691), .ZN(n7679) );
  NAND2X0 U6924 ( .IN1(n7692), .IN2(n7693), .QN(n7676) );
  AO222X1 U6925 ( .IN1(n7694), .IN2(n7695), .IN3(n7696), .IN4(n7697), .IN5(
        n7698), .IN6(n7699), .Q(n7693) );
  AO222X1 U6926 ( .IN1(n7700), .IN2(n7701), .IN3(n7702), .IN4(n7703), .IN5(
        n7704), .IN6(n7705), .Q(n7697) );
  AO22X1 U6927 ( .IN1(n7706), .IN2(n7707), .IN3(n7708), .IN4(n7709), .Q(n7702)
         );
  MUX21X1 U6928 ( .IN1(n7710), .IN2(n7711), .S(n7712), .Q(n7707) );
  AO222X1 U6929 ( .IN1(n7713), .IN2(n7714), .IN3(n7715), .IN4(n7716), .IN5(
        n7717), .IN6(n7718), .Q(n7710) );
  AO222X1 U6930 ( .IN1(n7719), .IN2(n7720), .IN3(n7721), .IN4(n7722), .IN5(
        n7723), .IN6(n7724), .Q(n7715) );
  AO221X1 U6931 ( .IN1(n7725), .IN2(n7726), .IN3(n7727), .IN4(n7728), .IN5(
        n7729), .Q(n7721) );
  AO222X1 U6932 ( .IN1(n7730), .IN2(n7731), .IN3(n7732), .IN4(n7733), .IN5(
        n7734), .IN6(n7735), .Q(n7729) );
  AO222X1 U6933 ( .IN1(n7736), .IN2(n7737), .IN3(n7738), .IN4(n7739), .IN5(
        n7740), .IN6(n7741), .Q(n7734) );
  AO222X1 U6934 ( .IN1(n7742), .IN2(n7743), .IN3(n7744), .IN4(n7745), .IN5(
        n7746), .IN6(n7747), .Q(n7738) );
  OAI222X1 U6935 ( .IN1(n7748), .IN2(n7749), .IN3(n7750), .IN4(n7751), .IN5(
        n7752), .IN6(n7753), .QN(n7744) );
  OA222X1 U6936 ( .IN1(n7754), .IN2(n7755), .IN3(n7756), .IN4(n7757), .IN5(
        n7758), .IN6(n7759), .Q(n7750) );
  OA222X1 U6937 ( .IN1(n7760), .IN2(n7761), .IN3(n7762), .IN4(n7664), .IN5(
        n7763), .IN6(n7764), .Q(n7756) );
  OA22X1 U6938 ( .IN1(n4485), .IN2(n7765), .IN3(n4484), .IN4(n7766), .Q(n7762)
         );
  OA21X1 U6939 ( .IN1(n7767), .IN2(n7768), .IN3(n5695), .Q(n7673) );
  AND3X1 U6940 ( .IN1(n7399), .IN2(n7521), .IN3(N4809), .Q(n7768) );
  AND3X1 U6941 ( .IN1(n7769), .IN2(n7770), .IN3(N4845), .Q(n7767) );
  AO22X1 U6942 ( .IN1(n3723), .IN2(n7771), .IN3(n7400), .IN4(n7772), .Q(n7561)
         );
  NAND4X0 U6943 ( .IN1(n7773), .IN2(n7774), .IN3(n7775), .IN4(n7776), .QN(
        n7772) );
  NAND3X0 U6944 ( .IN1(n7777), .IN2(n3720), .IN3(N1767), .QN(n7776) );
  NAND3X0 U6945 ( .IN1(n7576), .IN2(n7526), .IN3(N4710), .QN(n7775) );
  NAND2X0 U6946 ( .IN1(N4776), .IN2(n7778), .QN(n7774) );
  MUX21X1 U6947 ( .IN1(n7779), .IN2(n7780), .S(n3721), .Q(n7773) );
  NAND2X0 U6948 ( .IN1(N4677), .IN2(n7399), .QN(n7780) );
  OA22X1 U6949 ( .IN1(n7395), .IN2(n7781), .IN3(n7782), .IN4(n7573), .Q(n7779)
         );
  INVX0 U6950 ( .INP(N4513), .ZN(n7573) );
  AO221X1 U6951 ( .IN1(N4743), .IN2(n7783), .IN3(n7784), .IN4(n7785), .IN5(
        n7786), .Q(n7771) );
  MUX21X1 U6952 ( .IN1(n7787), .IN2(n7788), .S(n3719), .Q(n7786) );
  NOR2X0 U6953 ( .IN1(n7789), .IN2(n7782), .QN(n7788) );
  AOI22X1 U6954 ( .IN1(n7545), .IN2(N1767), .IN3(n3721), .IN4(N4611), .QN(
        n7789) );
  AND2X1 U6955 ( .IN1(N5292), .IN2(n5696), .Q(n7787) );
  AO222X1 U6956 ( .IN1(N1767), .IN2(n7576), .IN3(n506), .IN4(n7545), .IN5(n393), .IN6(n3720), .Q(n7785) );
  OAI22X1 U6957 ( .IN1(n7394), .IN2(n7457), .IN3(n7458), .IN4(n3720), .QN(
        n7783) );
  OA22X1 U6958 ( .IN1(n7790), .IN2(n7791), .IN3(n7792), .IN4(n7521), .Q(n7559)
         );
  OA221X1 U6959 ( .IN1(n7793), .IN2(n7530), .IN3(n7781), .IN4(n7794), .IN5(
        n7795), .Q(n7792) );
  NAND4X0 U6960 ( .IN1(N4915), .IN2(n7769), .IN3(n7777), .IN4(n7450), .QN(
        n7795) );
  NAND2X0 U6961 ( .IN1(n7778), .IN2(n3721), .QN(n7794) );
  INVX0 U6962 ( .INP(N4546), .ZN(n7781) );
  AOI22X1 U6963 ( .IN1(n7452), .IN2(n506), .IN3(n7513), .IN4(n393), .QN(n7793)
         );
  INVX0 U6964 ( .INP(N1767), .ZN(n7791) );
  OA221X1 U6965 ( .IN1(n3719), .IN2(n7796), .IN3(n7797), .IN4(n7798), .IN5(
        n7509), .Q(n7790) );
  NAND2X0 U6966 ( .IN1(n7770), .IN2(n7401), .QN(n7509) );
  NAND2X0 U6967 ( .IN1(n7450), .IN2(n5695), .QN(n7798) );
  AOI22X1 U6968 ( .IN1(n3721), .IN2(n7778), .IN3(n7799), .IN4(n7576), .QN(
        n7796) );
  INVX0 U6969 ( .INP(n7800), .ZN(n7778) );
  NAND3X0 U6970 ( .IN1(n7399), .IN2(n7401), .IN3(n506), .QN(n7558) );
  NAND2X0 U6971 ( .IN1(N5194), .IN2(n7801), .QN(n7557) );
  AO222X1 U6972 ( .IN1(n7802), .IN2(n538), .IN3(n7803), .IN4(n425), .IN5(n9122), .IN6(n7804), .Q(n4140) );
  AO222X1 U6973 ( .IN1(n7802), .IN2(n537), .IN3(n424), .IN4(n7803), .IN5(n9121), .IN6(n7804), .Q(n4139) );
  AO222X1 U6974 ( .IN1(n7092), .IN2(n537), .IN3(n7805), .IN4(n424), .IN5(n9120), .IN6(n7093), .Q(n4138) );
  AO222X1 U6975 ( .IN1(n7802), .IN2(n536), .IN3(n423), .IN4(n7803), .IN5(n9119), .IN6(n7804), .Q(n4137) );
  AO222X1 U6976 ( .IN1(n7092), .IN2(n536), .IN3(n423), .IN4(n7805), .IN5(n9118), .IN6(n7093), .Q(n4136) );
  AO222X1 U6977 ( .IN1(n7802), .IN2(n535), .IN3(n422), .IN4(n7803), .IN5(n9117), .IN6(n7804), .Q(n4135) );
  AO222X1 U6978 ( .IN1(n7092), .IN2(n535), .IN3(n422), .IN4(n7805), .IN5(n9116), .IN6(n7093), .Q(n4134) );
  AO222X1 U6979 ( .IN1(n7802), .IN2(n534), .IN3(n421), .IN4(n7803), .IN5(n9115), .IN6(n7804), .Q(n4133) );
  AO222X1 U6980 ( .IN1(n7092), .IN2(n534), .IN3(n421), .IN4(n7805), .IN5(n9114), .IN6(n7093), .Q(n4132) );
  AO222X1 U6981 ( .IN1(n7802), .IN2(n533), .IN3(n420), .IN4(n7803), .IN5(n9113), .IN6(n7804), .Q(n4131) );
  AO222X1 U6982 ( .IN1(n7092), .IN2(n533), .IN3(n420), .IN4(n7805), .IN5(n9112), .IN6(n7093), .Q(n4130) );
  AO222X1 U6983 ( .IN1(n7802), .IN2(n532), .IN3(n419), .IN4(n7803), .IN5(n9111), .IN6(n7804), .Q(n4129) );
  AO222X1 U6984 ( .IN1(n7092), .IN2(n532), .IN3(n419), .IN4(n7805), .IN5(n9110), .IN6(n7093), .Q(n4128) );
  AO222X1 U6985 ( .IN1(n7802), .IN2(n531), .IN3(n418), .IN4(n7803), .IN5(n9109), .IN6(n7804), .Q(n4127) );
  AO222X1 U6986 ( .IN1(n7092), .IN2(n531), .IN3(n418), .IN4(n7805), .IN5(n9108), .IN6(n7093), .Q(n4126) );
  AO222X1 U6987 ( .IN1(n7802), .IN2(n530), .IN3(n417), .IN4(n7803), .IN5(n9107), .IN6(n7804), .Q(n4125) );
  AO222X1 U6988 ( .IN1(n7092), .IN2(n530), .IN3(n417), .IN4(n7805), .IN5(n9106), .IN6(n7093), .Q(n4124) );
  AO222X1 U6989 ( .IN1(n7802), .IN2(n529), .IN3(n416), .IN4(n7803), .IN5(n9105), .IN6(n7804), .Q(n4123) );
  AO222X1 U6990 ( .IN1(n7092), .IN2(n529), .IN3(n416), .IN4(n7805), .IN5(n9104), .IN6(n7093), .Q(n4122) );
  AO222X1 U6991 ( .IN1(n7802), .IN2(n528), .IN3(n415), .IN4(n7803), .IN5(n9103), .IN6(n7804), .Q(n4121) );
  AO222X1 U6992 ( .IN1(n7092), .IN2(n528), .IN3(n415), .IN4(n7805), .IN5(n9102), .IN6(n7093), .Q(n4120) );
  AO222X1 U6993 ( .IN1(n7802), .IN2(n527), .IN3(n414), .IN4(n7803), .IN5(n9101), .IN6(n7804), .Q(n4119) );
  AO222X1 U6994 ( .IN1(n7092), .IN2(n527), .IN3(n414), .IN4(n7805), .IN5(n9100), .IN6(n7093), .Q(n4118) );
  AO222X1 U6995 ( .IN1(n7802), .IN2(n526), .IN3(n413), .IN4(n7803), .IN5(n9099), .IN6(n7804), .Q(n4117) );
  AO222X1 U6996 ( .IN1(n7092), .IN2(n526), .IN3(n413), .IN4(n7805), .IN5(n9098), .IN6(n7093), .Q(n4116) );
  AO222X1 U6997 ( .IN1(n7802), .IN2(n525), .IN3(n412), .IN4(n7803), .IN5(n9097), .IN6(n7804), .Q(n4115) );
  AO222X1 U6998 ( .IN1(n7092), .IN2(n525), .IN3(n412), .IN4(n7805), .IN5(n9096), .IN6(n7093), .Q(n4114) );
  AO222X1 U6999 ( .IN1(n7802), .IN2(n524), .IN3(n411), .IN4(n7803), .IN5(n9095), .IN6(n7804), .Q(n4113) );
  AO222X1 U7000 ( .IN1(n7092), .IN2(n524), .IN3(n411), .IN4(n7805), .IN5(n9094), .IN6(n7093), .Q(n4112) );
  AO222X1 U7001 ( .IN1(n7802), .IN2(n523), .IN3(n410), .IN4(n7803), .IN5(n9093), .IN6(n7804), .Q(n4111) );
  AO222X1 U7002 ( .IN1(n7092), .IN2(n523), .IN3(n410), .IN4(n7805), .IN5(n9092), .IN6(n7093), .Q(n4110) );
  AO222X1 U7003 ( .IN1(n7802), .IN2(n522), .IN3(n409), .IN4(n7803), .IN5(n9091), .IN6(n7804), .Q(n4109) );
  AO222X1 U7004 ( .IN1(n7092), .IN2(n522), .IN3(n409), .IN4(n7805), .IN5(n9090), .IN6(n7093), .Q(n4108) );
  AO222X1 U7005 ( .IN1(n7802), .IN2(n521), .IN3(n408), .IN4(n7803), .IN5(n9089), .IN6(n7804), .Q(n4107) );
  AO222X1 U7006 ( .IN1(n7092), .IN2(n521), .IN3(n408), .IN4(n7805), .IN5(n9088), .IN6(n7093), .Q(n4106) );
  AO222X1 U7007 ( .IN1(n7802), .IN2(n520), .IN3(n407), .IN4(n7803), .IN5(n9087), .IN6(n7804), .Q(n4105) );
  AO222X1 U7008 ( .IN1(n7092), .IN2(n520), .IN3(n407), .IN4(n7805), .IN5(n9086), .IN6(n7093), .Q(n4104) );
  AO222X1 U7009 ( .IN1(n7802), .IN2(n519), .IN3(n406), .IN4(n7803), .IN5(n9085), .IN6(n7804), .Q(n4103) );
  AO222X1 U7010 ( .IN1(n7092), .IN2(n519), .IN3(n406), .IN4(n7805), .IN5(n9084), .IN6(n7093), .Q(n4102) );
  AO222X1 U7011 ( .IN1(n7802), .IN2(n518), .IN3(n405), .IN4(n7803), .IN5(n9083), .IN6(n7804), .Q(n4101) );
  AO222X1 U7012 ( .IN1(n7092), .IN2(n518), .IN3(n405), .IN4(n7805), .IN5(n9082), .IN6(n7093), .Q(n4100) );
  AO222X1 U7013 ( .IN1(n7802), .IN2(n517), .IN3(n404), .IN4(n7803), .IN5(n9081), .IN6(n7804), .Q(n4099) );
  AO222X1 U7014 ( .IN1(n7092), .IN2(n517), .IN3(n404), .IN4(n7805), .IN5(n9080), .IN6(n7093), .Q(n4098) );
  AO222X1 U7015 ( .IN1(n7802), .IN2(n516), .IN3(n403), .IN4(n7803), .IN5(n9079), .IN6(n7804), .Q(n4097) );
  AO222X1 U7016 ( .IN1(n7092), .IN2(n516), .IN3(n403), .IN4(n7805), .IN5(n9078), .IN6(n7093), .Q(n4096) );
  AO222X1 U7017 ( .IN1(n7802), .IN2(n515), .IN3(n402), .IN4(n7803), .IN5(n9077), .IN6(n7804), .Q(n4095) );
  AO222X1 U7018 ( .IN1(n7092), .IN2(n515), .IN3(n402), .IN4(n7805), .IN5(n9076), .IN6(n7093), .Q(n4094) );
  AO222X1 U7019 ( .IN1(n7802), .IN2(n514), .IN3(n401), .IN4(n7803), .IN5(n9075), .IN6(n7804), .Q(n4093) );
  AO222X1 U7020 ( .IN1(n7092), .IN2(n514), .IN3(n401), .IN4(n7805), .IN5(n9074), .IN6(n7093), .Q(n4092) );
  AO222X1 U7021 ( .IN1(n7802), .IN2(n513), .IN3(n400), .IN4(n7803), .IN5(n9073), .IN6(n7804), .Q(n4091) );
  AO222X1 U7022 ( .IN1(n7092), .IN2(n513), .IN3(n400), .IN4(n7805), .IN5(n9072), .IN6(n7093), .Q(n4090) );
  AO222X1 U7023 ( .IN1(n7802), .IN2(n512), .IN3(n399), .IN4(n7803), .IN5(n9071), .IN6(n7804), .Q(n4089) );
  AO222X1 U7024 ( .IN1(n7092), .IN2(n512), .IN3(n399), .IN4(n7805), .IN5(n9070), .IN6(n7093), .Q(n4088) );
  AO222X1 U7025 ( .IN1(n7802), .IN2(n511), .IN3(n398), .IN4(n7803), .IN5(n9069), .IN6(n7804), .Q(n4087) );
  AO222X1 U7026 ( .IN1(n7092), .IN2(n511), .IN3(n398), .IN4(n7805), .IN5(n9068), .IN6(n7093), .Q(n4086) );
  AO222X1 U7027 ( .IN1(n7802), .IN2(n510), .IN3(n397), .IN4(n7803), .IN5(n9067), .IN6(n7804), .Q(n4085) );
  AO222X1 U7028 ( .IN1(n7092), .IN2(n510), .IN3(n397), .IN4(n7805), .IN5(n9066), .IN6(n7093), .Q(n4084) );
  AO222X1 U7029 ( .IN1(n7802), .IN2(n509), .IN3(n396), .IN4(n7803), .IN5(n9065), .IN6(n7804), .Q(n4083) );
  AO222X1 U7030 ( .IN1(n7092), .IN2(n509), .IN3(n396), .IN4(n7805), .IN5(n9064), .IN6(n7093), .Q(n4082) );
  AO222X1 U7031 ( .IN1(n7802), .IN2(n508), .IN3(n395), .IN4(n7803), .IN5(n9063), .IN6(n7804), .Q(n4081) );
  AO222X1 U7032 ( .IN1(n7092), .IN2(n508), .IN3(n395), .IN4(n7805), .IN5(n9062), .IN6(n7093), .Q(n4080) );
  AO222X1 U7033 ( .IN1(n7802), .IN2(n507), .IN3(n394), .IN4(n7803), .IN5(n9061), .IN6(n7804), .Q(n4079) );
  AOI21X1 U7034 ( .IN1(n7806), .IN2(n7807), .IN3(n7804), .QN(n7803) );
  NAND2X0 U7035 ( .IN1(n3716), .IN2(\r1720/A[3] ), .QN(n7807) );
  NOR2X0 U7036 ( .IN1(n7804), .IN2(n7577), .QN(n7802) );
  NAND2X0 U7037 ( .IN1(n4419), .IN2(reset_n), .QN(n7804) );
  AOI21X1 U7038 ( .IN1(n7808), .IN2(n7809), .IN3(n9191), .QN(n4419) );
  NAND4X0 U7039 ( .IN1(n7401), .IN2(n7810), .IN3(n7521), .IN4(n5695), .QN(
        n7809) );
  AO21X1 U7040 ( .IN1(\r1720/A[3] ), .IN2(n7811), .IN3(n7399), .Q(n7810) );
  NAND2X0 U7041 ( .IN1(n7812), .IN2(n7526), .QN(n7808) );
  AO22X1 U7042 ( .IN1(n7524), .IN2(n7401), .IN3(n7813), .IN4(n7555), .Q(n7812)
         );
  NOR2X0 U7043 ( .IN1(n3719), .IN2(n7457), .QN(n7813) );
  MUX21X1 U7044 ( .IN1(IF_PC[31]), .IN2(N466), .S(reset_n), .Q(n4078) );
  MUX21X1 U7045 ( .IN1(IF_PC[0]), .IN2(N435), .S(reset_n), .Q(n4077) );
  MUX21X1 U7046 ( .IN1(IF_PC[1]), .IN2(N436), .S(reset_n), .Q(n4076) );
  MUX21X1 U7047 ( .IN1(IF_PC[2]), .IN2(N437), .S(reset_n), .Q(n4075) );
  MUX21X1 U7048 ( .IN1(IF_PC[3]), .IN2(N438), .S(reset_n), .Q(n4074) );
  MUX21X1 U7049 ( .IN1(IF_PC[4]), .IN2(N439), .S(reset_n), .Q(n4073) );
  MUX21X1 U7050 ( .IN1(IF_PC[5]), .IN2(N440), .S(reset_n), .Q(n4072) );
  MUX21X1 U7051 ( .IN1(IF_PC[6]), .IN2(N441), .S(reset_n), .Q(n4071) );
  MUX21X1 U7052 ( .IN1(IF_PC[7]), .IN2(N442), .S(reset_n), .Q(n4070) );
  MUX21X1 U7053 ( .IN1(IF_PC[8]), .IN2(N443), .S(reset_n), .Q(n4069) );
  MUX21X1 U7054 ( .IN1(IF_PC[9]), .IN2(N444), .S(reset_n), .Q(n4068) );
  MUX21X1 U7055 ( .IN1(IF_PC[10]), .IN2(N445), .S(reset_n), .Q(n4067) );
  MUX21X1 U7056 ( .IN1(IF_PC[11]), .IN2(N446), .S(reset_n), .Q(n4066) );
  MUX21X1 U7057 ( .IN1(IF_PC[12]), .IN2(N447), .S(reset_n), .Q(n4065) );
  MUX21X1 U7058 ( .IN1(IF_PC[13]), .IN2(N448), .S(reset_n), .Q(n4064) );
  MUX21X1 U7059 ( .IN1(IF_PC[14]), .IN2(N449), .S(reset_n), .Q(n4063) );
  MUX21X1 U7060 ( .IN1(IF_PC[15]), .IN2(N450), .S(reset_n), .Q(n4062) );
  MUX21X1 U7061 ( .IN1(IF_PC[16]), .IN2(N451), .S(reset_n), .Q(n4061) );
  MUX21X1 U7062 ( .IN1(IF_PC[17]), .IN2(N452), .S(reset_n), .Q(n4060) );
  MUX21X1 U7063 ( .IN1(IF_PC[18]), .IN2(N453), .S(reset_n), .Q(n4059) );
  MUX21X1 U7064 ( .IN1(IF_PC[19]), .IN2(N454), .S(reset_n), .Q(n4058) );
  MUX21X1 U7065 ( .IN1(IF_PC[20]), .IN2(N455), .S(reset_n), .Q(n4057) );
  MUX21X1 U7066 ( .IN1(IF_PC[21]), .IN2(N456), .S(reset_n), .Q(n4056) );
  MUX21X1 U7067 ( .IN1(IF_PC[22]), .IN2(N457), .S(reset_n), .Q(n4055) );
  MUX21X1 U7068 ( .IN1(IF_PC[23]), .IN2(N458), .S(reset_n), .Q(n4054) );
  MUX21X1 U7069 ( .IN1(IF_PC[24]), .IN2(N459), .S(reset_n), .Q(n4053) );
  MUX21X1 U7070 ( .IN1(IF_PC[25]), .IN2(N460), .S(reset_n), .Q(n4052) );
  MUX21X1 U7071 ( .IN1(IF_PC[26]), .IN2(N461), .S(reset_n), .Q(n4051) );
  MUX21X1 U7072 ( .IN1(IF_PC[27]), .IN2(N462), .S(reset_n), .Q(n4050) );
  MUX21X1 U7073 ( .IN1(IF_PC[28]), .IN2(N463), .S(reset_n), .Q(n4049) );
  MUX21X1 U7074 ( .IN1(IF_PC[29]), .IN2(N464), .S(reset_n), .Q(n4048) );
  MUX21X1 U7075 ( .IN1(IF_PC[30]), .IN2(N465), .S(reset_n), .Q(n4047) );
  AO221X1 U7076 ( .IN1(n7814), .IN2(N5622), .IN3(n7815), .IN4(n9156), .IN5(
        n7816), .Q(n4046) );
  AO22X1 U7077 ( .IN1(n9060), .IN2(n7817), .IN3(n7818), .IN4(n7263), .Q(n7816)
         );
  AO221X1 U7078 ( .IN1(n7814), .IN2(N5623), .IN3(n7815), .IN4(n9155), .IN5(
        n7819), .Q(n4045) );
  AO22X1 U7079 ( .IN1(n9059), .IN2(n7817), .IN3(n7818), .IN4(n7262), .Q(n7819)
         );
  AO221X1 U7080 ( .IN1(n7814), .IN2(N5624), .IN3(n7815), .IN4(n9154), .IN5(
        n7820), .Q(n4044) );
  AO22X1 U7081 ( .IN1(n9058), .IN2(n7817), .IN3(n7818), .IN4(n7261), .Q(n7820)
         );
  AO221X1 U7082 ( .IN1(n7814), .IN2(N5625), .IN3(n7815), .IN4(n9153), .IN5(
        n7821), .Q(n4043) );
  AO22X1 U7083 ( .IN1(n9057), .IN2(n7817), .IN3(n7818), .IN4(n7260), .Q(n7821)
         );
  AO221X1 U7084 ( .IN1(n7814), .IN2(N5626), .IN3(n7815), .IN4(n9152), .IN5(
        n7822), .Q(n4042) );
  AO22X1 U7085 ( .IN1(n9056), .IN2(n7817), .IN3(n7818), .IN4(n7259), .Q(n7822)
         );
  AO221X1 U7086 ( .IN1(n7814), .IN2(N5627), .IN3(n7815), .IN4(n9151), .IN5(
        n7823), .Q(n4041) );
  AO22X1 U7087 ( .IN1(n9055), .IN2(n7817), .IN3(n7818), .IN4(n7258), .Q(n7823)
         );
  AO221X1 U7088 ( .IN1(n7814), .IN2(N5628), .IN3(n7815), .IN4(n9150), .IN5(
        n7824), .Q(n4040) );
  AO22X1 U7089 ( .IN1(n9054), .IN2(n7817), .IN3(n7818), .IN4(n7257), .Q(n7824)
         );
  AO221X1 U7090 ( .IN1(n7814), .IN2(N5629), .IN3(n7815), .IN4(n9149), .IN5(
        n7825), .Q(n4039) );
  AO22X1 U7091 ( .IN1(n9053), .IN2(n7817), .IN3(n7818), .IN4(n7256), .Q(n7825)
         );
  AO221X1 U7092 ( .IN1(n7814), .IN2(N5630), .IN3(n7815), .IN4(n9148), .IN5(
        n7826), .Q(n4038) );
  AO22X1 U7093 ( .IN1(n9052), .IN2(n7817), .IN3(n7818), .IN4(n7255), .Q(n7826)
         );
  AO221X1 U7094 ( .IN1(n7814), .IN2(N5631), .IN3(n7815), .IN4(n9147), .IN5(
        n7827), .Q(n4037) );
  AO22X1 U7095 ( .IN1(n9051), .IN2(n7817), .IN3(n7818), .IN4(n7254), .Q(n7827)
         );
  AO221X1 U7096 ( .IN1(n7814), .IN2(N5632), .IN3(n7815), .IN4(n9146), .IN5(
        n7828), .Q(n4036) );
  AO22X1 U7097 ( .IN1(n9050), .IN2(n7817), .IN3(n7818), .IN4(n7253), .Q(n7828)
         );
  AO221X1 U7098 ( .IN1(n7814), .IN2(N5633), .IN3(n7815), .IN4(n9145), .IN5(
        n7829), .Q(n4035) );
  AO22X1 U7099 ( .IN1(n9049), .IN2(n7817), .IN3(n7818), .IN4(n7252), .Q(n7829)
         );
  AO221X1 U7100 ( .IN1(n7814), .IN2(N5634), .IN3(n7815), .IN4(n9144), .IN5(
        n7830), .Q(n4034) );
  AO22X1 U7101 ( .IN1(n9048), .IN2(n7817), .IN3(n7818), .IN4(n7251), .Q(n7830)
         );
  AO221X1 U7102 ( .IN1(n7814), .IN2(N5635), .IN3(n7815), .IN4(n9143), .IN5(
        n7831), .Q(n4033) );
  AO22X1 U7103 ( .IN1(n9047), .IN2(n7817), .IN3(n7818), .IN4(n7250), .Q(n7831)
         );
  AO221X1 U7104 ( .IN1(n7814), .IN2(N5636), .IN3(n7815), .IN4(n9142), .IN5(
        n7832), .Q(n4032) );
  AO22X1 U7105 ( .IN1(n9046), .IN2(n7817), .IN3(n7818), .IN4(n7249), .Q(n7832)
         );
  AO221X1 U7106 ( .IN1(n7814), .IN2(N5637), .IN3(n7815), .IN4(n9141), .IN5(
        n7833), .Q(n4031) );
  AO22X1 U7107 ( .IN1(n9045), .IN2(n7817), .IN3(n7818), .IN4(n7248), .Q(n7833)
         );
  AO221X1 U7108 ( .IN1(n7814), .IN2(N5638), .IN3(n7815), .IN4(n9140), .IN5(
        n7834), .Q(n4030) );
  AO22X1 U7109 ( .IN1(n9044), .IN2(n7817), .IN3(n7818), .IN4(n7247), .Q(n7834)
         );
  AO221X1 U7110 ( .IN1(n7814), .IN2(N5639), .IN3(n7815), .IN4(n9139), .IN5(
        n7835), .Q(n4029) );
  AO22X1 U7111 ( .IN1(n9043), .IN2(n7817), .IN3(n7818), .IN4(n7246), .Q(n7835)
         );
  AO221X1 U7112 ( .IN1(n7814), .IN2(N5640), .IN3(n7815), .IN4(n9138), .IN5(
        n7836), .Q(n4028) );
  AO22X1 U7113 ( .IN1(n9042), .IN2(n7817), .IN3(n7818), .IN4(n7245), .Q(n7836)
         );
  AO221X1 U7114 ( .IN1(n7814), .IN2(N5641), .IN3(n7815), .IN4(n9137), .IN5(
        n7837), .Q(n4027) );
  AO22X1 U7115 ( .IN1(n9041), .IN2(n7817), .IN3(n7818), .IN4(n7244), .Q(n7837)
         );
  AO221X1 U7116 ( .IN1(n7814), .IN2(N5642), .IN3(n7815), .IN4(n9136), .IN5(
        n7838), .Q(n4026) );
  AO22X1 U7117 ( .IN1(n9040), .IN2(n7817), .IN3(n7818), .IN4(n7243), .Q(n7838)
         );
  AO221X1 U7118 ( .IN1(n7814), .IN2(N5643), .IN3(n7815), .IN4(n9135), .IN5(
        n7839), .Q(n4025) );
  AO22X1 U7119 ( .IN1(n9039), .IN2(n7817), .IN3(n7818), .IN4(n7242), .Q(n7839)
         );
  AO221X1 U7120 ( .IN1(n7814), .IN2(N5644), .IN3(n7815), .IN4(n9134), .IN5(
        n7840), .Q(n4024) );
  AO22X1 U7121 ( .IN1(n9038), .IN2(n7817), .IN3(n7818), .IN4(n7241), .Q(n7840)
         );
  AO221X1 U7122 ( .IN1(n7814), .IN2(N5645), .IN3(n7815), .IN4(n9133), .IN5(
        n7841), .Q(n4023) );
  AO22X1 U7123 ( .IN1(n9037), .IN2(n7817), .IN3(n7818), .IN4(n7240), .Q(n7841)
         );
  AO221X1 U7124 ( .IN1(n7814), .IN2(N5646), .IN3(n7815), .IN4(n9132), .IN5(
        n7842), .Q(n4022) );
  AO22X1 U7125 ( .IN1(n9036), .IN2(n7817), .IN3(n7818), .IN4(n7239), .Q(n7842)
         );
  AO221X1 U7126 ( .IN1(n7814), .IN2(N5647), .IN3(n7815), .IN4(n9131), .IN5(
        n7843), .Q(n4021) );
  AO22X1 U7127 ( .IN1(n9035), .IN2(n7817), .IN3(n7818), .IN4(n7238), .Q(n7843)
         );
  AO221X1 U7128 ( .IN1(n7814), .IN2(N5648), .IN3(n7815), .IN4(n9130), .IN5(
        n7844), .Q(n4020) );
  AO22X1 U7129 ( .IN1(n9034), .IN2(n7817), .IN3(n7818), .IN4(n7237), .Q(n7844)
         );
  AO221X1 U7130 ( .IN1(n7814), .IN2(N5649), .IN3(n7815), .IN4(n9129), .IN5(
        n7845), .Q(n4019) );
  AO22X1 U7131 ( .IN1(n9033), .IN2(n7817), .IN3(n7818), .IN4(n7236), .Q(n7845)
         );
  AO221X1 U7132 ( .IN1(n7814), .IN2(N5650), .IN3(n7815), .IN4(n9128), .IN5(
        n7846), .Q(n4018) );
  AO22X1 U7133 ( .IN1(n9032), .IN2(n7817), .IN3(n7818), .IN4(n7235), .Q(n7846)
         );
  AO221X1 U7134 ( .IN1(n7814), .IN2(N5651), .IN3(n7815), .IN4(n9127), .IN5(
        n7847), .Q(n4017) );
  AO22X1 U7135 ( .IN1(n9031), .IN2(n7817), .IN3(n7818), .IN4(n7234), .Q(n7847)
         );
  AO221X1 U7136 ( .IN1(n7814), .IN2(N5652), .IN3(n7815), .IN4(n9126), .IN5(
        n7848), .Q(n4016) );
  AO22X1 U7137 ( .IN1(n9030), .IN2(n7817), .IN3(n7818), .IN4(n7233), .Q(n7848)
         );
  AND2X1 U7138 ( .IN1(n7849), .IN2(n7441), .Q(n7815) );
  AND2X1 U7139 ( .IN1(n7849), .IN2(n7850), .Q(n7814) );
  AO222X1 U7140 ( .IN1(n7849), .IN2(n7101), .IN3(n7818), .IN4(n7232), .IN5(
        n9029), .IN6(n7817), .Q(n4015) );
  AND3X1 U7141 ( .IN1(n7527), .IN2(n7801), .IN3(n7851), .Q(n7818) );
  INVX0 U7142 ( .INP(n7852), .ZN(n7801) );
  MUX21X1 U7143 ( .IN1(N5653), .IN2(n9125), .S(n7441), .Q(n7101) );
  INVX0 U7144 ( .INP(n7850), .ZN(n7441) );
  NAND3X0 U7145 ( .IN1(n7449), .IN2(n7853), .IN3(n7854), .QN(n7850) );
  OA222X1 U7146 ( .IN1(n7545), .IN2(n7499), .IN3(n7401), .IN4(n7855), .IN5(
        n7856), .IN6(n7531), .Q(n7854) );
  NOR2X0 U7147 ( .IN1(n7526), .IN2(n7811), .QN(n7856) );
  INVX0 U7148 ( .INP(n7857), .ZN(n7811) );
  MUX21X1 U7149 ( .IN1(n7858), .IN2(n7859), .S(n9167), .Q(n7857) );
  MUX21X1 U7150 ( .IN1(n7860), .IN2(n7861), .S(n9168), .Q(n7859) );
  NOR2X0 U7151 ( .IN1(n9190), .IN2(n7862), .QN(n7861) );
  XNOR2X1 U7152 ( .IN1(n9166), .IN2(n7863), .Q(n7862) );
  MUX21X1 U7153 ( .IN1(n7864), .IN2(n7865), .S(n9123), .Q(n7860) );
  NAND2X0 U7154 ( .IN1(n9166), .IN2(n7866), .QN(n7865) );
  OR2X1 U7155 ( .IN1(n7866), .IN2(n9166), .Q(n7864) );
  MUX21X1 U7156 ( .IN1(n4486), .IN2(n7863), .S(n9190), .Q(n7866) );
  XOR2X1 U7157 ( .IN1(n9169), .IN2(n9124), .Q(n7863) );
  XNOR2X1 U7158 ( .IN1(n9166), .IN2(n7867), .Q(n7858) );
  MUX41X1 U7159 ( .IN1(n9123), .IN3(n9173), .IN2(n9124), .IN4(n9169), .S0(
        n9168), .S1(n9190), .Q(n7867) );
  AND2X1 U7160 ( .IN1(n7868), .IN2(n7869), .Q(n7855) );
  NAND2X0 U7161 ( .IN1(n7451), .IN2(n7550), .QN(n7853) );
  OA21X1 U7162 ( .IN1(n3716), .IN2(n3719), .IN3(n7870), .Q(n7449) );
  AND2X1 U7163 ( .IN1(n7851), .IN2(n7871), .Q(n7849) );
  NAND3X0 U7164 ( .IN1(n7538), .IN2(n7470), .IN3(n7872), .QN(n7871) );
  OA221X1 U7165 ( .IN1(n7868), .IN2(n7471), .IN3(n7527), .IN4(n7852), .IN5(
        n7873), .Q(n7872) );
  NAND3X0 U7166 ( .IN1(n7513), .IN2(n7874), .IN3(n7450), .QN(n7873) );
  NAND2X0 U7167 ( .IN1(n7524), .IN2(n3720), .QN(n7852) );
  INVX0 U7168 ( .INP(n7540), .ZN(n7524) );
  NAND2X0 U7169 ( .IN1(n7577), .IN2(n7521), .QN(n7540) );
  INVX0 U7170 ( .INP(n7531), .ZN(n7577) );
  NOR2X0 U7171 ( .IN1(n7875), .IN2(n7271), .QN(n7527) );
  OA221X1 U7172 ( .IN1(n7876), .IN2(n7512), .IN3(n7877), .IN4(n7508), .IN5(
        n7878), .Q(n7470) );
  OA21X1 U7173 ( .IN1(n3716), .IN2(n7544), .IN3(n7542), .Q(n7878) );
  AOI21X1 U7174 ( .IN1(n7879), .IN2(n7521), .IN3(n7880), .QN(n7542) );
  NOR4X0 U7175 ( .IN1(n3719), .IN2(n3716), .IN3(n7881), .IN4(n5753), .QN(n7880) );
  OA21X1 U7176 ( .IN1(n3720), .IN2(n3723), .IN3(n7806), .Q(n7881) );
  NAND2X0 U7177 ( .IN1(n7882), .IN2(n7883), .QN(n7879) );
  NAND3X0 U7178 ( .IN1(n3716), .IN2(n7497), .IN3(n7513), .QN(n7883) );
  NAND3X0 U7179 ( .IN1(n7401), .IN2(n3723), .IN3(n7777), .QN(n7882) );
  NAND3X0 U7180 ( .IN1(n3719), .IN2(n5753), .IN3(n7452), .QN(n7544) );
  OA222X1 U7181 ( .IN1(n7884), .IN2(n7550), .IN3(n3721), .IN4(n7868), .IN5(
        n7885), .IN6(n7806), .Q(n7877) );
  INVX0 U7182 ( .INP(n7497), .ZN(n7885) );
  NAND2X0 U7183 ( .IN1(n7457), .IN2(n7530), .QN(n7497) );
  NAND2X0 U7184 ( .IN1(\r1720/A[3] ), .IN2(n5695), .QN(n7868) );
  AOI22X1 U7185 ( .IN1(n7447), .IN2(n7500), .IN3(n7511), .IN4(n7451), .QN(
        n7876) );
  NOR2X0 U7186 ( .IN1(n7884), .IN2(n3719), .QN(n7500) );
  AOI22X1 U7187 ( .IN1(n7532), .IN2(n7452), .IN3(n7886), .IN4(n7513), .QN(
        n7538) );
  NOR2X0 U7188 ( .IN1(n5753), .IN2(n7870), .QN(n7886) );
  NOR2X0 U7189 ( .IN1(n5695), .IN2(\r1720/A[3] ), .QN(n7452) );
  INVX0 U7190 ( .INP(n7471), .ZN(n7532) );
  INVX0 U7191 ( .INP(n7817), .ZN(n7851) );
  NAND2X0 U7192 ( .IN1(n7114), .IN2(n7442), .QN(n7817) );
  NAND4X0 U7193 ( .IN1(n7471), .IN2(n7579), .IN3(n7887), .IN4(n7888), .QN(
        n7442) );
  OA22X1 U7194 ( .IN1(n3721), .IN2(n7889), .IN3(n7450), .IN4(n7549), .Q(n7888)
         );
  AO21X1 U7195 ( .IN1(n7508), .IN2(n7447), .IN3(n7512), .Q(n7887) );
  NAND2X0 U7196 ( .IN1(n7511), .IN2(n7457), .QN(n7471) );
  INVX0 U7197 ( .INP(n7870), .ZN(n7511) );
  AO222X1 U7198 ( .IN1(n7092), .IN2(n507), .IN3(n394), .IN4(n7805), .IN5(n9028), .IN6(n7093), .Q(n4014) );
  NOR2X0 U7199 ( .IN1(n7093), .IN2(n5695), .QN(n7805) );
  NOR2X0 U7200 ( .IN1(n7093), .IN2(n3723), .QN(n7092) );
  NAND4X0 U7201 ( .IN1(n7890), .IN2(n7401), .IN3(n7114), .IN4(n7556), .QN(
        n7093) );
  INVX0 U7202 ( .INP(n7097), .ZN(n7114) );
  NAND2X0 U7203 ( .IN1(reset_n), .IN2(n5701), .QN(n7097) );
  INVX0 U7204 ( .INP(n7530), .ZN(n7401) );
  NAND2X0 U7205 ( .IN1(n3721), .IN2(n3720), .QN(n7530) );
  MUX21X1 U7206 ( .IN1(n7399), .IN2(n7770), .S(n3723), .Q(n7890) );
  MUX21X1 U7207 ( .IN1(n7891), .IN2(\R[7][31] ), .S(n7892), .Q(n4013) );
  MUX21X1 U7208 ( .IN1(n7893), .IN2(\R[7][30] ), .S(n7892), .Q(n4012) );
  MUX21X1 U7209 ( .IN1(n7894), .IN2(\R[7][29] ), .S(n7892), .Q(n4011) );
  MUX21X1 U7210 ( .IN1(n7895), .IN2(\R[7][28] ), .S(n7892), .Q(n4010) );
  MUX21X1 U7211 ( .IN1(n7896), .IN2(\R[7][27] ), .S(n7892), .Q(n4009) );
  MUX21X1 U7212 ( .IN1(n7897), .IN2(\R[7][26] ), .S(n7892), .Q(n4008) );
  MUX21X1 U7213 ( .IN1(n7898), .IN2(\R[7][25] ), .S(n7892), .Q(n4007) );
  MUX21X1 U7214 ( .IN1(n7899), .IN2(\R[7][24] ), .S(n7892), .Q(n4006) );
  MUX21X1 U7215 ( .IN1(n7900), .IN2(\R[7][23] ), .S(n7892), .Q(n4005) );
  MUX21X1 U7216 ( .IN1(n7901), .IN2(\R[7][22] ), .S(n7892), .Q(n4004) );
  MUX21X1 U7217 ( .IN1(n7902), .IN2(\R[7][21] ), .S(n7892), .Q(n4003) );
  MUX21X1 U7218 ( .IN1(n7903), .IN2(\R[7][20] ), .S(n7892), .Q(n4002) );
  MUX21X1 U7219 ( .IN1(n7904), .IN2(\R[7][19] ), .S(n7892), .Q(n4001) );
  MUX21X1 U7220 ( .IN1(n7905), .IN2(\R[7][18] ), .S(n7892), .Q(n4000) );
  MUX21X1 U7221 ( .IN1(n7906), .IN2(\R[7][17] ), .S(n7892), .Q(n3999) );
  MUX21X1 U7222 ( .IN1(n7907), .IN2(\R[7][16] ), .S(n7892), .Q(n3998) );
  MUX21X1 U7223 ( .IN1(n7908), .IN2(\R[7][15] ), .S(n7892), .Q(n3997) );
  MUX21X1 U7224 ( .IN1(n7909), .IN2(\R[7][14] ), .S(n7892), .Q(n3996) );
  MUX21X1 U7225 ( .IN1(n7910), .IN2(\R[7][13] ), .S(n7892), .Q(n3995) );
  MUX21X1 U7226 ( .IN1(n7911), .IN2(\R[7][12] ), .S(n7892), .Q(n3994) );
  MUX21X1 U7227 ( .IN1(n7912), .IN2(\R[7][11] ), .S(n7892), .Q(n3993) );
  MUX21X1 U7228 ( .IN1(n7913), .IN2(\R[7][10] ), .S(n7892), .Q(n3992) );
  MUX21X1 U7229 ( .IN1(n7914), .IN2(\R[7][9] ), .S(n7892), .Q(n3991) );
  MUX21X1 U7230 ( .IN1(n7915), .IN2(\R[7][8] ), .S(n7892), .Q(n3990) );
  MUX21X1 U7231 ( .IN1(n7916), .IN2(\R[7][7] ), .S(n7892), .Q(n3989) );
  MUX21X1 U7232 ( .IN1(n7917), .IN2(\R[7][6] ), .S(n7892), .Q(n3988) );
  MUX21X1 U7233 ( .IN1(n7918), .IN2(\R[7][5] ), .S(n7892), .Q(n3987) );
  MUX21X1 U7234 ( .IN1(n7919), .IN2(\R[7][4] ), .S(n7892), .Q(n3986) );
  MUX21X1 U7235 ( .IN1(n7920), .IN2(\R[7][3] ), .S(n7892), .Q(n3985) );
  MUX21X1 U7236 ( .IN1(n7921), .IN2(\R[7][2] ), .S(n7892), .Q(n3984) );
  MUX21X1 U7237 ( .IN1(n7922), .IN2(\R[7][1] ), .S(n7892), .Q(n3983) );
  MUX21X1 U7238 ( .IN1(n7923), .IN2(\R[7][0] ), .S(n7892), .Q(n3982) );
  AND2X1 U7239 ( .IN1(n7924), .IN2(n7925), .Q(n7892) );
  NAND3X0 U7240 ( .IN1(n7926), .IN2(n7927), .IN3(n7928), .QN(n7925) );
  NAND3X0 U7241 ( .IN1(n9161), .IN2(n9162), .IN3(n7929), .QN(n7924) );
  MUX21X1 U7242 ( .IN1(n7891), .IN2(\R[6][31] ), .S(n7930), .Q(n3981) );
  MUX21X1 U7243 ( .IN1(n7893), .IN2(\R[6][30] ), .S(n7930), .Q(n3980) );
  MUX21X1 U7244 ( .IN1(n7894), .IN2(\R[6][29] ), .S(n7930), .Q(n3979) );
  MUX21X1 U7245 ( .IN1(n7895), .IN2(\R[6][28] ), .S(n7930), .Q(n3978) );
  MUX21X1 U7246 ( .IN1(n7896), .IN2(\R[6][27] ), .S(n7930), .Q(n3977) );
  MUX21X1 U7247 ( .IN1(n7897), .IN2(\R[6][26] ), .S(n7930), .Q(n3976) );
  MUX21X1 U7248 ( .IN1(n7898), .IN2(\R[6][25] ), .S(n7930), .Q(n3975) );
  MUX21X1 U7249 ( .IN1(n7899), .IN2(\R[6][24] ), .S(n7930), .Q(n3974) );
  MUX21X1 U7250 ( .IN1(n7900), .IN2(\R[6][23] ), .S(n7930), .Q(n3973) );
  MUX21X1 U7251 ( .IN1(n7901), .IN2(\R[6][22] ), .S(n7930), .Q(n3972) );
  MUX21X1 U7252 ( .IN1(n7902), .IN2(\R[6][21] ), .S(n7930), .Q(n3971) );
  MUX21X1 U7253 ( .IN1(n7903), .IN2(\R[6][20] ), .S(n7930), .Q(n3970) );
  MUX21X1 U7254 ( .IN1(n7904), .IN2(\R[6][19] ), .S(n7930), .Q(n3969) );
  MUX21X1 U7255 ( .IN1(n7905), .IN2(\R[6][18] ), .S(n7930), .Q(n3968) );
  MUX21X1 U7256 ( .IN1(n7906), .IN2(\R[6][17] ), .S(n7930), .Q(n3967) );
  MUX21X1 U7257 ( .IN1(n7907), .IN2(\R[6][16] ), .S(n7930), .Q(n3966) );
  MUX21X1 U7258 ( .IN1(n7908), .IN2(\R[6][15] ), .S(n7930), .Q(n3965) );
  MUX21X1 U7259 ( .IN1(n7909), .IN2(\R[6][14] ), .S(n7930), .Q(n3964) );
  MUX21X1 U7260 ( .IN1(n7910), .IN2(\R[6][13] ), .S(n7930), .Q(n3963) );
  MUX21X1 U7261 ( .IN1(n7911), .IN2(\R[6][12] ), .S(n7930), .Q(n3962) );
  MUX21X1 U7262 ( .IN1(n7912), .IN2(\R[6][11] ), .S(n7930), .Q(n3961) );
  MUX21X1 U7263 ( .IN1(n7913), .IN2(\R[6][10] ), .S(n7930), .Q(n3960) );
  MUX21X1 U7264 ( .IN1(n7914), .IN2(\R[6][9] ), .S(n7930), .Q(n3959) );
  MUX21X1 U7265 ( .IN1(n7915), .IN2(\R[6][8] ), .S(n7930), .Q(n3958) );
  MUX21X1 U7266 ( .IN1(n7916), .IN2(\R[6][7] ), .S(n7930), .Q(n3957) );
  MUX21X1 U7267 ( .IN1(n7917), .IN2(\R[6][6] ), .S(n7930), .Q(n3956) );
  MUX21X1 U7268 ( .IN1(n7918), .IN2(\R[6][5] ), .S(n7930), .Q(n3955) );
  MUX21X1 U7269 ( .IN1(n7919), .IN2(\R[6][4] ), .S(n7930), .Q(n3954) );
  MUX21X1 U7270 ( .IN1(n7920), .IN2(\R[6][3] ), .S(n7930), .Q(n3953) );
  MUX21X1 U7271 ( .IN1(n7921), .IN2(\R[6][2] ), .S(n7930), .Q(n3952) );
  MUX21X1 U7272 ( .IN1(n7922), .IN2(\R[6][1] ), .S(n7930), .Q(n3951) );
  MUX21X1 U7273 ( .IN1(n7923), .IN2(\R[6][0] ), .S(n7930), .Q(n3950) );
  AND2X1 U7274 ( .IN1(n7931), .IN2(n7932), .Q(n7930) );
  NAND3X0 U7275 ( .IN1(n7928), .IN2(n7926), .IN3(n7933), .QN(n7932) );
  NAND3X0 U7276 ( .IN1(n9161), .IN2(n5704), .IN3(n7929), .QN(n7931) );
  MUX21X1 U7277 ( .IN1(n7891), .IN2(\R[5][31] ), .S(n7934), .Q(n3949) );
  MUX21X1 U7278 ( .IN1(n7893), .IN2(\R[5][30] ), .S(n7934), .Q(n3948) );
  MUX21X1 U7279 ( .IN1(n7894), .IN2(\R[5][29] ), .S(n7934), .Q(n3947) );
  MUX21X1 U7280 ( .IN1(n7895), .IN2(\R[5][28] ), .S(n7934), .Q(n3946) );
  MUX21X1 U7281 ( .IN1(n7896), .IN2(\R[5][27] ), .S(n7934), .Q(n3945) );
  MUX21X1 U7282 ( .IN1(n7897), .IN2(\R[5][26] ), .S(n7934), .Q(n3944) );
  MUX21X1 U7283 ( .IN1(n7898), .IN2(\R[5][25] ), .S(n7934), .Q(n3943) );
  MUX21X1 U7284 ( .IN1(n7899), .IN2(\R[5][24] ), .S(n7934), .Q(n3942) );
  MUX21X1 U7285 ( .IN1(n7900), .IN2(\R[5][23] ), .S(n7934), .Q(n3941) );
  MUX21X1 U7286 ( .IN1(n7901), .IN2(\R[5][22] ), .S(n7934), .Q(n3940) );
  MUX21X1 U7287 ( .IN1(n7902), .IN2(\R[5][21] ), .S(n7934), .Q(n3939) );
  MUX21X1 U7288 ( .IN1(n7903), .IN2(\R[5][20] ), .S(n7934), .Q(n3938) );
  MUX21X1 U7289 ( .IN1(n7904), .IN2(\R[5][19] ), .S(n7934), .Q(n3937) );
  MUX21X1 U7290 ( .IN1(n7905), .IN2(\R[5][18] ), .S(n7934), .Q(n3936) );
  MUX21X1 U7291 ( .IN1(n7906), .IN2(\R[5][17] ), .S(n7934), .Q(n3935) );
  MUX21X1 U7292 ( .IN1(n7907), .IN2(\R[5][16] ), .S(n7934), .Q(n3934) );
  MUX21X1 U7293 ( .IN1(n7908), .IN2(\R[5][15] ), .S(n7934), .Q(n3933) );
  MUX21X1 U7294 ( .IN1(n7909), .IN2(\R[5][14] ), .S(n7934), .Q(n3932) );
  MUX21X1 U7295 ( .IN1(n7910), .IN2(\R[5][13] ), .S(n7934), .Q(n3931) );
  MUX21X1 U7296 ( .IN1(n7911), .IN2(\R[5][12] ), .S(n7934), .Q(n3930) );
  MUX21X1 U7297 ( .IN1(n7912), .IN2(\R[5][11] ), .S(n7934), .Q(n3929) );
  MUX21X1 U7298 ( .IN1(n7913), .IN2(\R[5][10] ), .S(n7934), .Q(n3928) );
  MUX21X1 U7299 ( .IN1(n7914), .IN2(\R[5][9] ), .S(n7934), .Q(n3927) );
  MUX21X1 U7300 ( .IN1(n7915), .IN2(\R[5][8] ), .S(n7934), .Q(n3926) );
  MUX21X1 U7301 ( .IN1(n7916), .IN2(\R[5][7] ), .S(n7934), .Q(n3925) );
  MUX21X1 U7302 ( .IN1(n7917), .IN2(\R[5][6] ), .S(n7934), .Q(n3924) );
  MUX21X1 U7303 ( .IN1(n7918), .IN2(\R[5][5] ), .S(n7934), .Q(n3923) );
  MUX21X1 U7304 ( .IN1(n7919), .IN2(\R[5][4] ), .S(n7934), .Q(n3922) );
  MUX21X1 U7305 ( .IN1(n7920), .IN2(\R[5][3] ), .S(n7934), .Q(n3921) );
  MUX21X1 U7306 ( .IN1(n7921), .IN2(\R[5][2] ), .S(n7934), .Q(n3920) );
  MUX21X1 U7307 ( .IN1(n7922), .IN2(\R[5][1] ), .S(n7934), .Q(n3919) );
  MUX21X1 U7308 ( .IN1(n7923), .IN2(\R[5][0] ), .S(n7934), .Q(n3918) );
  AND2X1 U7309 ( .IN1(n7935), .IN2(n7936), .Q(n7934) );
  NAND3X0 U7310 ( .IN1(n7926), .IN2(n7927), .IN3(n7937), .QN(n7936) );
  NAND3X0 U7311 ( .IN1(n9162), .IN2(n5691), .IN3(n7929), .QN(n7935) );
  MUX21X1 U7312 ( .IN1(n7891), .IN2(\R[4][31] ), .S(n7938), .Q(n3917) );
  MUX21X1 U7313 ( .IN1(n7893), .IN2(\R[4][30] ), .S(n7938), .Q(n3916) );
  MUX21X1 U7314 ( .IN1(n7894), .IN2(\R[4][29] ), .S(n7938), .Q(n3915) );
  MUX21X1 U7315 ( .IN1(n7895), .IN2(\R[4][28] ), .S(n7938), .Q(n3914) );
  MUX21X1 U7316 ( .IN1(n7896), .IN2(\R[4][27] ), .S(n7938), .Q(n3913) );
  MUX21X1 U7317 ( .IN1(n7897), .IN2(\R[4][26] ), .S(n7938), .Q(n3912) );
  MUX21X1 U7318 ( .IN1(n7898), .IN2(\R[4][25] ), .S(n7938), .Q(n3911) );
  MUX21X1 U7319 ( .IN1(n7899), .IN2(\R[4][24] ), .S(n7938), .Q(n3910) );
  MUX21X1 U7320 ( .IN1(n7900), .IN2(\R[4][23] ), .S(n7938), .Q(n3909) );
  MUX21X1 U7321 ( .IN1(n7901), .IN2(\R[4][22] ), .S(n7938), .Q(n3908) );
  MUX21X1 U7322 ( .IN1(n7902), .IN2(\R[4][21] ), .S(n7938), .Q(n3907) );
  MUX21X1 U7323 ( .IN1(n7903), .IN2(\R[4][20] ), .S(n7938), .Q(n3906) );
  MUX21X1 U7324 ( .IN1(n7904), .IN2(\R[4][19] ), .S(n7938), .Q(n3905) );
  MUX21X1 U7325 ( .IN1(n7905), .IN2(\R[4][18] ), .S(n7938), .Q(n3904) );
  MUX21X1 U7326 ( .IN1(n7906), .IN2(\R[4][17] ), .S(n7938), .Q(n3903) );
  MUX21X1 U7327 ( .IN1(n7907), .IN2(\R[4][16] ), .S(n7938), .Q(n3902) );
  MUX21X1 U7328 ( .IN1(n7908), .IN2(\R[4][15] ), .S(n7938), .Q(n3901) );
  MUX21X1 U7329 ( .IN1(n7909), .IN2(\R[4][14] ), .S(n7938), .Q(n3900) );
  MUX21X1 U7330 ( .IN1(n7910), .IN2(\R[4][13] ), .S(n7938), .Q(n3899) );
  MUX21X1 U7331 ( .IN1(n7911), .IN2(\R[4][12] ), .S(n7938), .Q(n3898) );
  MUX21X1 U7332 ( .IN1(n7912), .IN2(\R[4][11] ), .S(n7938), .Q(n3897) );
  MUX21X1 U7333 ( .IN1(n7913), .IN2(\R[4][10] ), .S(n7938), .Q(n3896) );
  MUX21X1 U7334 ( .IN1(n7914), .IN2(\R[4][9] ), .S(n7938), .Q(n3895) );
  MUX21X1 U7335 ( .IN1(n7915), .IN2(\R[4][8] ), .S(n7938), .Q(n3894) );
  MUX21X1 U7336 ( .IN1(n7916), .IN2(\R[4][7] ), .S(n7938), .Q(n3893) );
  MUX21X1 U7337 ( .IN1(n7917), .IN2(\R[4][6] ), .S(n7938), .Q(n3892) );
  MUX21X1 U7338 ( .IN1(n7918), .IN2(\R[4][5] ), .S(n7938), .Q(n3891) );
  MUX21X1 U7339 ( .IN1(n7919), .IN2(\R[4][4] ), .S(n7938), .Q(n3890) );
  MUX21X1 U7340 ( .IN1(n7920), .IN2(\R[4][3] ), .S(n7938), .Q(n3889) );
  MUX21X1 U7341 ( .IN1(n7921), .IN2(\R[4][2] ), .S(n7938), .Q(n3888) );
  MUX21X1 U7342 ( .IN1(n7922), .IN2(\R[4][1] ), .S(n7938), .Q(n3887) );
  MUX21X1 U7343 ( .IN1(n7923), .IN2(\R[4][0] ), .S(n7938), .Q(n3886) );
  AND2X1 U7344 ( .IN1(n7939), .IN2(n7940), .Q(n7938) );
  NAND3X0 U7345 ( .IN1(n7933), .IN2(n7926), .IN3(n7937), .QN(n7940) );
  NAND3X0 U7346 ( .IN1(n5704), .IN2(n5691), .IN3(n7929), .QN(n7939) );
  AND2X1 U7347 ( .IN1(n9160), .IN2(n7941), .Q(n7929) );
  MUX21X1 U7348 ( .IN1(n7891), .IN2(\R[3][31] ), .S(n7942), .Q(n3885) );
  MUX21X1 U7349 ( .IN1(n7893), .IN2(\R[3][30] ), .S(n7942), .Q(n3884) );
  MUX21X1 U7350 ( .IN1(n7894), .IN2(\R[3][29] ), .S(n7942), .Q(n3883) );
  MUX21X1 U7351 ( .IN1(n7895), .IN2(\R[3][28] ), .S(n7942), .Q(n3882) );
  MUX21X1 U7352 ( .IN1(n7896), .IN2(\R[3][27] ), .S(n7942), .Q(n3881) );
  MUX21X1 U7353 ( .IN1(n7897), .IN2(\R[3][26] ), .S(n7942), .Q(n3880) );
  MUX21X1 U7354 ( .IN1(n7898), .IN2(\R[3][25] ), .S(n7942), .Q(n3879) );
  MUX21X1 U7355 ( .IN1(n7899), .IN2(\R[3][24] ), .S(n7942), .Q(n3878) );
  MUX21X1 U7356 ( .IN1(n7900), .IN2(\R[3][23] ), .S(n7942), .Q(n3877) );
  MUX21X1 U7357 ( .IN1(n7901), .IN2(\R[3][22] ), .S(n7942), .Q(n3876) );
  MUX21X1 U7358 ( .IN1(n7902), .IN2(\R[3][21] ), .S(n7942), .Q(n3875) );
  MUX21X1 U7359 ( .IN1(n7903), .IN2(\R[3][20] ), .S(n7942), .Q(n3874) );
  MUX21X1 U7360 ( .IN1(n7904), .IN2(\R[3][19] ), .S(n7942), .Q(n3873) );
  MUX21X1 U7361 ( .IN1(n7905), .IN2(\R[3][18] ), .S(n7942), .Q(n3872) );
  MUX21X1 U7362 ( .IN1(n7906), .IN2(\R[3][17] ), .S(n7942), .Q(n3871) );
  MUX21X1 U7363 ( .IN1(n7907), .IN2(\R[3][16] ), .S(n7942), .Q(n3870) );
  MUX21X1 U7364 ( .IN1(n7908), .IN2(\R[3][15] ), .S(n7942), .Q(n3869) );
  MUX21X1 U7365 ( .IN1(n7909), .IN2(\R[3][14] ), .S(n7942), .Q(n3868) );
  MUX21X1 U7366 ( .IN1(n7910), .IN2(\R[3][13] ), .S(n7942), .Q(n3867) );
  MUX21X1 U7367 ( .IN1(n7911), .IN2(\R[3][12] ), .S(n7942), .Q(n3866) );
  MUX21X1 U7368 ( .IN1(n7912), .IN2(\R[3][11] ), .S(n7942), .Q(n3865) );
  MUX21X1 U7369 ( .IN1(n7913), .IN2(\R[3][10] ), .S(n7942), .Q(n3864) );
  MUX21X1 U7370 ( .IN1(n7914), .IN2(\R[3][9] ), .S(n7942), .Q(n3863) );
  MUX21X1 U7371 ( .IN1(n7915), .IN2(\R[3][8] ), .S(n7942), .Q(n3862) );
  MUX21X1 U7372 ( .IN1(n7916), .IN2(\R[3][7] ), .S(n7942), .Q(n3861) );
  MUX21X1 U7373 ( .IN1(n7917), .IN2(\R[3][6] ), .S(n7942), .Q(n3860) );
  MUX21X1 U7374 ( .IN1(n7918), .IN2(\R[3][5] ), .S(n7942), .Q(n3859) );
  MUX21X1 U7375 ( .IN1(n7919), .IN2(\R[3][4] ), .S(n7942), .Q(n3858) );
  MUX21X1 U7376 ( .IN1(n7920), .IN2(\R[3][3] ), .S(n7942), .Q(n3857) );
  MUX21X1 U7377 ( .IN1(n7921), .IN2(\R[3][2] ), .S(n7942), .Q(n3856) );
  MUX21X1 U7378 ( .IN1(n7922), .IN2(\R[3][1] ), .S(n7942), .Q(n3855) );
  MUX21X1 U7379 ( .IN1(n7923), .IN2(\R[3][0] ), .S(n7942), .Q(n3854) );
  AND2X1 U7380 ( .IN1(n7943), .IN2(n7944), .Q(n7942) );
  NAND3X0 U7381 ( .IN1(n7928), .IN2(n7927), .IN3(n7945), .QN(n7944) );
  NAND3X0 U7382 ( .IN1(n9161), .IN2(n9162), .IN3(n7946), .QN(n7943) );
  MUX21X1 U7383 ( .IN1(n7891), .IN2(\R[2][31] ), .S(n7947), .Q(n3853) );
  MUX21X1 U7384 ( .IN1(n7893), .IN2(\R[2][30] ), .S(n7947), .Q(n3852) );
  MUX21X1 U7385 ( .IN1(n7894), .IN2(\R[2][29] ), .S(n7947), .Q(n3851) );
  MUX21X1 U7386 ( .IN1(n7895), .IN2(\R[2][28] ), .S(n7947), .Q(n3850) );
  MUX21X1 U7387 ( .IN1(n7896), .IN2(\R[2][27] ), .S(n7947), .Q(n3849) );
  MUX21X1 U7388 ( .IN1(n7897), .IN2(\R[2][26] ), .S(n7947), .Q(n3848) );
  MUX21X1 U7389 ( .IN1(n7898), .IN2(\R[2][25] ), .S(n7947), .Q(n3847) );
  MUX21X1 U7390 ( .IN1(n7899), .IN2(\R[2][24] ), .S(n7947), .Q(n3846) );
  MUX21X1 U7391 ( .IN1(n7900), .IN2(\R[2][23] ), .S(n7947), .Q(n3845) );
  MUX21X1 U7392 ( .IN1(n7901), .IN2(\R[2][22] ), .S(n7947), .Q(n3844) );
  MUX21X1 U7393 ( .IN1(n7902), .IN2(\R[2][21] ), .S(n7947), .Q(n3843) );
  MUX21X1 U7394 ( .IN1(n7903), .IN2(\R[2][20] ), .S(n7947), .Q(n3842) );
  MUX21X1 U7395 ( .IN1(n7904), .IN2(\R[2][19] ), .S(n7947), .Q(n3841) );
  MUX21X1 U7396 ( .IN1(n7905), .IN2(\R[2][18] ), .S(n7947), .Q(n3840) );
  MUX21X1 U7397 ( .IN1(n7906), .IN2(\R[2][17] ), .S(n7947), .Q(n3839) );
  MUX21X1 U7398 ( .IN1(n7907), .IN2(\R[2][16] ), .S(n7947), .Q(n3838) );
  MUX21X1 U7399 ( .IN1(n7908), .IN2(\R[2][15] ), .S(n7947), .Q(n3837) );
  MUX21X1 U7400 ( .IN1(n7909), .IN2(\R[2][14] ), .S(n7947), .Q(n3836) );
  MUX21X1 U7401 ( .IN1(n7910), .IN2(\R[2][13] ), .S(n7947), .Q(n3835) );
  MUX21X1 U7402 ( .IN1(n7911), .IN2(\R[2][12] ), .S(n7947), .Q(n3834) );
  MUX21X1 U7403 ( .IN1(n7912), .IN2(\R[2][11] ), .S(n7947), .Q(n3833) );
  MUX21X1 U7404 ( .IN1(n7913), .IN2(\R[2][10] ), .S(n7947), .Q(n3832) );
  MUX21X1 U7405 ( .IN1(n7914), .IN2(\R[2][9] ), .S(n7947), .Q(n3831) );
  MUX21X1 U7406 ( .IN1(n7915), .IN2(\R[2][8] ), .S(n7947), .Q(n3830) );
  MUX21X1 U7407 ( .IN1(n7916), .IN2(\R[2][7] ), .S(n7947), .Q(n3829) );
  MUX21X1 U7408 ( .IN1(n7917), .IN2(\R[2][6] ), .S(n7947), .Q(n3828) );
  MUX21X1 U7409 ( .IN1(n7918), .IN2(\R[2][5] ), .S(n7947), .Q(n3827) );
  MUX21X1 U7410 ( .IN1(n7919), .IN2(\R[2][4] ), .S(n7947), .Q(n3826) );
  MUX21X1 U7411 ( .IN1(n7920), .IN2(\R[2][3] ), .S(n7947), .Q(n3825) );
  MUX21X1 U7412 ( .IN1(n7921), .IN2(\R[2][2] ), .S(n7947), .Q(n3824) );
  MUX21X1 U7413 ( .IN1(n7922), .IN2(\R[2][1] ), .S(n7947), .Q(n3823) );
  MUX21X1 U7414 ( .IN1(n7923), .IN2(\R[2][0] ), .S(n7947), .Q(n3822) );
  AND2X1 U7415 ( .IN1(n7948), .IN2(n7949), .Q(n7947) );
  NAND3X0 U7416 ( .IN1(n7933), .IN2(n7928), .IN3(n7945), .QN(n7949) );
  AND2X1 U7417 ( .IN1(n7950), .IN2(n7951), .Q(n7928) );
  NAND3X0 U7418 ( .IN1(n9161), .IN2(n5704), .IN3(n7946), .QN(n7948) );
  MUX21X1 U7419 ( .IN1(n7891), .IN2(\R[1][31] ), .S(n7952), .Q(n3821) );
  MUX21X1 U7420 ( .IN1(n7893), .IN2(\R[1][30] ), .S(n7952), .Q(n3820) );
  MUX21X1 U7421 ( .IN1(n7894), .IN2(\R[1][29] ), .S(n7952), .Q(n3819) );
  MUX21X1 U7422 ( .IN1(n7895), .IN2(\R[1][28] ), .S(n7952), .Q(n3818) );
  MUX21X1 U7423 ( .IN1(n7896), .IN2(\R[1][27] ), .S(n7952), .Q(n3817) );
  MUX21X1 U7424 ( .IN1(n7897), .IN2(\R[1][26] ), .S(n7952), .Q(n3816) );
  MUX21X1 U7425 ( .IN1(n7898), .IN2(\R[1][25] ), .S(n7952), .Q(n3815) );
  MUX21X1 U7426 ( .IN1(n7899), .IN2(\R[1][24] ), .S(n7952), .Q(n3814) );
  MUX21X1 U7427 ( .IN1(n7900), .IN2(\R[1][23] ), .S(n7952), .Q(n3813) );
  MUX21X1 U7428 ( .IN1(n7901), .IN2(\R[1][22] ), .S(n7952), .Q(n3812) );
  MUX21X1 U7429 ( .IN1(n7902), .IN2(\R[1][21] ), .S(n7952), .Q(n3811) );
  MUX21X1 U7430 ( .IN1(n7903), .IN2(\R[1][20] ), .S(n7952), .Q(n3810) );
  MUX21X1 U7431 ( .IN1(n7904), .IN2(\R[1][19] ), .S(n7952), .Q(n3809) );
  MUX21X1 U7432 ( .IN1(n7905), .IN2(\R[1][18] ), .S(n7952), .Q(n3808) );
  MUX21X1 U7433 ( .IN1(n7906), .IN2(\R[1][17] ), .S(n7952), .Q(n3807) );
  MUX21X1 U7434 ( .IN1(n7907), .IN2(\R[1][16] ), .S(n7952), .Q(n3806) );
  MUX21X1 U7435 ( .IN1(n7908), .IN2(\R[1][15] ), .S(n7952), .Q(n3805) );
  MUX21X1 U7436 ( .IN1(n7909), .IN2(\R[1][14] ), .S(n7952), .Q(n3804) );
  MUX21X1 U7437 ( .IN1(n7910), .IN2(\R[1][13] ), .S(n7952), .Q(n3803) );
  MUX21X1 U7438 ( .IN1(n7911), .IN2(\R[1][12] ), .S(n7952), .Q(n3802) );
  MUX21X1 U7439 ( .IN1(n7912), .IN2(\R[1][11] ), .S(n7952), .Q(n3801) );
  MUX21X1 U7440 ( .IN1(n7913), .IN2(\R[1][10] ), .S(n7952), .Q(n3800) );
  MUX21X1 U7441 ( .IN1(n7914), .IN2(\R[1][9] ), .S(n7952), .Q(n3799) );
  MUX21X1 U7442 ( .IN1(n7915), .IN2(\R[1][8] ), .S(n7952), .Q(n3798) );
  MUX21X1 U7443 ( .IN1(n7916), .IN2(\R[1][7] ), .S(n7952), .Q(n3797) );
  MUX21X1 U7444 ( .IN1(n7917), .IN2(\R[1][6] ), .S(n7952), .Q(n3796) );
  MUX21X1 U7445 ( .IN1(n7918), .IN2(\R[1][5] ), .S(n7952), .Q(n3795) );
  MUX21X1 U7446 ( .IN1(n7919), .IN2(\R[1][4] ), .S(n7952), .Q(n3794) );
  MUX21X1 U7447 ( .IN1(n7920), .IN2(\R[1][3] ), .S(n7952), .Q(n3793) );
  MUX21X1 U7448 ( .IN1(n7921), .IN2(\R[1][2] ), .S(n7952), .Q(n3792) );
  MUX21X1 U7449 ( .IN1(n7922), .IN2(\R[1][1] ), .S(n7952), .Q(n3791) );
  MUX21X1 U7450 ( .IN1(n7923), .IN2(\R[1][0] ), .S(n7952), .Q(n3790) );
  AND2X1 U7451 ( .IN1(n7953), .IN2(n7954), .Q(n7952) );
  NAND3X0 U7452 ( .IN1(n7937), .IN2(n7927), .IN3(n7945), .QN(n7954) );
  INVX0 U7453 ( .INP(n7933), .ZN(n7927) );
  NAND3X0 U7454 ( .IN1(n9162), .IN2(n5691), .IN3(n7946), .QN(n7953) );
  MUX21X1 U7455 ( .IN1(n7891), .IN2(\R[0][31] ), .S(n7955), .Q(n3789) );
  AO221X1 U7456 ( .IN1(data[31]), .IN2(n7956), .IN3(n9029), .IN4(n7957), .IN5(
        n7958), .Q(n7891) );
  MUX21X1 U7457 ( .IN1(n7893), .IN2(\R[0][30] ), .S(n7955), .Q(n3788) );
  AO221X1 U7458 ( .IN1(data[30]), .IN2(n7956), .IN3(n9030), .IN4(n7957), .IN5(
        n7958), .Q(n7893) );
  MUX21X1 U7459 ( .IN1(n7894), .IN2(\R[0][29] ), .S(n7955), .Q(n3787) );
  AO221X1 U7460 ( .IN1(data[29]), .IN2(n7956), .IN3(n9031), .IN4(n7957), .IN5(
        n7958), .Q(n7894) );
  MUX21X1 U7461 ( .IN1(n7895), .IN2(\R[0][28] ), .S(n7955), .Q(n3786) );
  AO221X1 U7462 ( .IN1(data[28]), .IN2(n7956), .IN3(n9032), .IN4(n7957), .IN5(
        n7958), .Q(n7895) );
  MUX21X1 U7463 ( .IN1(n7896), .IN2(\R[0][27] ), .S(n7955), .Q(n3785) );
  AO221X1 U7464 ( .IN1(data[27]), .IN2(n7956), .IN3(n9033), .IN4(n7957), .IN5(
        n7958), .Q(n7896) );
  MUX21X1 U7465 ( .IN1(n7897), .IN2(\R[0][26] ), .S(n7955), .Q(n3784) );
  AO221X1 U7466 ( .IN1(data[26]), .IN2(n7956), .IN3(n9034), .IN4(n7957), .IN5(
        n7958), .Q(n7897) );
  MUX21X1 U7467 ( .IN1(n7898), .IN2(\R[0][25] ), .S(n7955), .Q(n3783) );
  AO221X1 U7468 ( .IN1(data[25]), .IN2(n7956), .IN3(n9035), .IN4(n7957), .IN5(
        n7958), .Q(n7898) );
  MUX21X1 U7469 ( .IN1(n7899), .IN2(\R[0][24] ), .S(n7955), .Q(n3782) );
  AO221X1 U7470 ( .IN1(data[24]), .IN2(n7956), .IN3(n9036), .IN4(n7957), .IN5(
        n7958), .Q(n7899) );
  MUX21X1 U7471 ( .IN1(n7900), .IN2(\R[0][23] ), .S(n7955), .Q(n3781) );
  AO221X1 U7472 ( .IN1(data[23]), .IN2(n7956), .IN3(n9037), .IN4(n7957), .IN5(
        n7958), .Q(n7900) );
  MUX21X1 U7473 ( .IN1(n7901), .IN2(\R[0][22] ), .S(n7955), .Q(n3780) );
  AO221X1 U7474 ( .IN1(data[22]), .IN2(n7956), .IN3(n9038), .IN4(n7957), .IN5(
        n7958), .Q(n7901) );
  MUX21X1 U7475 ( .IN1(n7902), .IN2(\R[0][21] ), .S(n7955), .Q(n3779) );
  AO221X1 U7476 ( .IN1(data[21]), .IN2(n7956), .IN3(n9039), .IN4(n7957), .IN5(
        n7958), .Q(n7902) );
  MUX21X1 U7477 ( .IN1(n7903), .IN2(\R[0][20] ), .S(n7955), .Q(n3778) );
  AO221X1 U7478 ( .IN1(data[20]), .IN2(n7956), .IN3(n9040), .IN4(n7957), .IN5(
        n7958), .Q(n7903) );
  MUX21X1 U7479 ( .IN1(n7904), .IN2(\R[0][19] ), .S(n7955), .Q(n3777) );
  AO221X1 U7480 ( .IN1(data[19]), .IN2(n7956), .IN3(n9041), .IN4(n7957), .IN5(
        n7958), .Q(n7904) );
  MUX21X1 U7481 ( .IN1(n7905), .IN2(\R[0][18] ), .S(n7955), .Q(n3776) );
  AO221X1 U7482 ( .IN1(data[18]), .IN2(n7956), .IN3(n9042), .IN4(n7957), .IN5(
        n7958), .Q(n7905) );
  MUX21X1 U7483 ( .IN1(n7906), .IN2(\R[0][17] ), .S(n7955), .Q(n3775) );
  AO221X1 U7484 ( .IN1(data[17]), .IN2(n7956), .IN3(n9043), .IN4(n7957), .IN5(
        n7958), .Q(n7906) );
  MUX21X1 U7485 ( .IN1(n7907), .IN2(\R[0][16] ), .S(n7955), .Q(n3774) );
  AO221X1 U7486 ( .IN1(data[16]), .IN2(n7956), .IN3(n9044), .IN4(n7957), .IN5(
        n7958), .Q(n7907) );
  NAND2X0 U7487 ( .IN1(n7959), .IN2(n7960), .QN(n7958) );
  NAND3X0 U7488 ( .IN1(n7961), .IN2(n9180), .IN3(data[15]), .QN(n7960) );
  NOR2X0 U7489 ( .IN1(n7962), .IN2(n7963), .QN(n7956) );
  INVX0 U7490 ( .INP(n7964), .ZN(n7963) );
  MUX21X1 U7491 ( .IN1(n7908), .IN2(\R[0][15] ), .S(n7955), .Q(n3773) );
  AO221X1 U7492 ( .IN1(data[15]), .IN2(n7965), .IN3(n9045), .IN4(n7957), .IN5(
        n7966), .Q(n7908) );
  MUX21X1 U7493 ( .IN1(n7909), .IN2(\R[0][14] ), .S(n7955), .Q(n3772) );
  AO221X1 U7494 ( .IN1(data[14]), .IN2(n7965), .IN3(n9046), .IN4(n7957), .IN5(
        n7966), .Q(n7909) );
  MUX21X1 U7495 ( .IN1(n7910), .IN2(\R[0][13] ), .S(n7955), .Q(n3771) );
  AO221X1 U7496 ( .IN1(data[13]), .IN2(n7965), .IN3(n9047), .IN4(n7957), .IN5(
        n7966), .Q(n7910) );
  MUX21X1 U7497 ( .IN1(n7911), .IN2(\R[0][12] ), .S(n7955), .Q(n3770) );
  AO221X1 U7498 ( .IN1(data[12]), .IN2(n7965), .IN3(n9048), .IN4(n7957), .IN5(
        n7966), .Q(n7911) );
  MUX21X1 U7499 ( .IN1(n7912), .IN2(\R[0][11] ), .S(n7955), .Q(n3769) );
  AO221X1 U7500 ( .IN1(data[11]), .IN2(n7965), .IN3(n9049), .IN4(n7957), .IN5(
        n7966), .Q(n7912) );
  MUX21X1 U7501 ( .IN1(n7913), .IN2(\R[0][10] ), .S(n7955), .Q(n3768) );
  AO221X1 U7502 ( .IN1(data[10]), .IN2(n7965), .IN3(n9050), .IN4(n7957), .IN5(
        n7966), .Q(n7913) );
  MUX21X1 U7503 ( .IN1(n7914), .IN2(\R[0][9] ), .S(n7955), .Q(n3767) );
  AO221X1 U7504 ( .IN1(data[9]), .IN2(n7965), .IN3(n9051), .IN4(n7957), .IN5(
        n7966), .Q(n7914) );
  MUX21X1 U7505 ( .IN1(n7915), .IN2(\R[0][8] ), .S(n7955), .Q(n3766) );
  AO221X1 U7506 ( .IN1(data[8]), .IN2(n7965), .IN3(n9052), .IN4(n7957), .IN5(
        n7966), .Q(n7915) );
  INVX0 U7507 ( .INP(n7959), .ZN(n7966) );
  NAND4X0 U7508 ( .IN1(data[7]), .IN2(n7961), .IN3(n9181), .IN4(n5708), .QN(
        n7959) );
  AO21X1 U7509 ( .IN1(n7967), .IN2(n7968), .IN3(n7950), .Q(n7965) );
  NAND2X0 U7510 ( .IN1(n7969), .IN2(n7962), .QN(n7968) );
  MUX21X1 U7511 ( .IN1(n7970), .IN2(n7971), .S(n9179), .Q(n7969) );
  NAND2X0 U7512 ( .IN1(n9180), .IN2(n9183), .QN(n7970) );
  MUX21X1 U7513 ( .IN1(n7916), .IN2(\R[0][7] ), .S(n7955), .Q(n3765) );
  AO22X1 U7514 ( .IN1(n9053), .IN2(n7957), .IN3(n7972), .IN4(data[7]), .Q(
        n7916) );
  MUX21X1 U7515 ( .IN1(n7917), .IN2(\R[0][6] ), .S(n7955), .Q(n3764) );
  AO22X1 U7516 ( .IN1(n9054), .IN2(n7957), .IN3(data[6]), .IN4(n7972), .Q(
        n7917) );
  MUX21X1 U7517 ( .IN1(n7918), .IN2(\R[0][5] ), .S(n7955), .Q(n3763) );
  AO22X1 U7518 ( .IN1(n9055), .IN2(n7957), .IN3(data[5]), .IN4(n7972), .Q(
        n7918) );
  MUX21X1 U7519 ( .IN1(n7919), .IN2(\R[0][4] ), .S(n7955), .Q(n3762) );
  AO22X1 U7520 ( .IN1(n9056), .IN2(n7957), .IN3(data[4]), .IN4(n7972), .Q(
        n7919) );
  MUX21X1 U7521 ( .IN1(n7920), .IN2(\R[0][3] ), .S(n7955), .Q(n3761) );
  AO22X1 U7522 ( .IN1(n9057), .IN2(n7957), .IN3(data[3]), .IN4(n7972), .Q(
        n7920) );
  MUX21X1 U7523 ( .IN1(n7921), .IN2(\R[0][2] ), .S(n7955), .Q(n3760) );
  AO22X1 U7524 ( .IN1(n9058), .IN2(n7957), .IN3(data[2]), .IN4(n7972), .Q(
        n7921) );
  MUX21X1 U7525 ( .IN1(n7922), .IN2(\R[0][1] ), .S(n7955), .Q(n3759) );
  AO22X1 U7526 ( .IN1(n9059), .IN2(n7957), .IN3(data[1]), .IN4(n7972), .Q(
        n7922) );
  MUX21X1 U7527 ( .IN1(n7923), .IN2(\R[0][0] ), .S(n7955), .Q(n3758) );
  AND2X1 U7528 ( .IN1(n7973), .IN2(n7974), .Q(n7955) );
  NAND3X0 U7529 ( .IN1(n7937), .IN2(n7933), .IN3(n7945), .QN(n7974) );
  INVX0 U7530 ( .INP(n7926), .ZN(n7945) );
  NAND4X0 U7531 ( .IN1(n5690), .IN2(n5687), .IN3(n5713), .IN4(n5694), .QN(
        n7926) );
  OA21X1 U7532 ( .IN1(n7975), .IN2(n9159), .IN3(n5687), .Q(n7933) );
  OA21X1 U7533 ( .IN1(n7976), .IN2(n9158), .IN3(n5690), .Q(n7975) );
  AOI21X1 U7534 ( .IN1(n5714), .IN2(n9176), .IN3(n9178), .QN(n7976) );
  NOR2X0 U7535 ( .IN1(n7951), .IN2(n7977), .QN(n7937) );
  INVX0 U7536 ( .INP(n7950), .ZN(n7977) );
  NOR4X0 U7537 ( .IN1(n7978), .IN2(n7962), .IN3(n5707), .IN4(n9181), .QN(n7950) );
  NAND3X0 U7538 ( .IN1(n5687), .IN2(n5713), .IN3(n7979), .QN(n7951) );
  NAND3X0 U7539 ( .IN1(n5690), .IN2(n5694), .IN3(n7980), .QN(n7979) );
  OR2X1 U7540 ( .IN1(n9177), .IN2(n9178), .Q(n7980) );
  NAND3X0 U7541 ( .IN1(n5704), .IN2(n5691), .IN3(n7946), .QN(n7973) );
  NOR2X0 U7542 ( .IN1(n7981), .IN2(n9160), .QN(n7946) );
  INVX0 U7543 ( .INP(n7941), .ZN(n7981) );
  AO21X1 U7544 ( .IN1(n7967), .IN2(n7982), .IN3(n7957), .Q(n7941) );
  NAND3X0 U7545 ( .IN1(n7983), .IN2(n7962), .IN3(n7971), .QN(n7982) );
  INVX0 U7546 ( .INP(n7961), .ZN(n7983) );
  AO22X1 U7547 ( .IN1(n9060), .IN2(n7957), .IN3(data[0]), .IN4(n7972), .Q(
        n7923) );
  AND3X1 U7548 ( .IN1(n7964), .IN2(n7984), .IN3(n7985), .Q(n7972) );
  OA22X1 U7549 ( .IN1(n7986), .IN2(n5707), .IN3(n5688), .IN4(n7987), .Q(n7985)
         );
  NOR2X0 U7550 ( .IN1(n5693), .IN2(n5688), .QN(n7986) );
  AO21X1 U7551 ( .IN1(n9182), .IN2(n5703), .IN3(n7967), .Q(n7964) );
  NOR2X0 U7552 ( .IN1(n5703), .IN2(n9182), .QN(n7967) );
  AO21X1 U7553 ( .IN1(n7988), .IN2(n5703), .IN3(n7989), .Q(n7957) );
  MUX21X1 U7554 ( .IN1(n7990), .IN2(n7991), .S(n9182), .Q(n7989) );
  NOR2X0 U7555 ( .IN1(n7992), .IN2(n5703), .QN(n7991) );
  MUX21X1 U7556 ( .IN1(n7962), .IN2(n7971), .S(n7993), .Q(n7992) );
  NOR2X0 U7557 ( .IN1(n9180), .IN2(n9179), .QN(n7993) );
  NAND2X0 U7558 ( .IN1(n9183), .IN2(n5710), .QN(n7962) );
  NOR2X0 U7559 ( .IN1(n7994), .IN2(n5688), .QN(n7990) );
  OA22X1 U7560 ( .IN1(n9180), .IN2(n7984), .IN3(n5703), .IN4(n7987), .Q(n7994)
         );
  AO221X1 U7561 ( .IN1(n7961), .IN2(n5708), .IN3(n7995), .IN4(n7978), .IN5(
        n7996), .Q(n7988) );
  MUX21X1 U7562 ( .IN1(n7997), .IN2(n7998), .S(n9182), .Q(n7996) );
  NOR2X0 U7563 ( .IN1(n7978), .IN2(n7971), .QN(n7998) );
  NAND2X0 U7564 ( .IN1(n9184), .IN2(n5693), .QN(n7971) );
  AO22X1 U7565 ( .IN1(n9180), .IN2(n5710), .IN3(n7987), .IN4(n5688), .Q(n7997)
         );
  NAND2X0 U7566 ( .IN1(n9180), .IN2(n9179), .QN(n7978) );
  INVX0 U7567 ( .INP(n7984), .ZN(n7995) );
  NAND2X0 U7568 ( .IN1(n5693), .IN2(n5710), .QN(n7984) );
  NOR2X0 U7569 ( .IN1(n7987), .IN2(n9179), .QN(n7961) );
  NAND2X0 U7570 ( .IN1(n9184), .IN2(n9183), .QN(n7987) );
  NAND2X0 U7571 ( .IN1(n3723), .IN2(n7870), .QN(n7999) );
  NOR2X0 U7572 ( .IN1(n3698), .IN2(n7782), .QN(\U3/U92/Z_9 ) );
  AO22X1 U7573 ( .IN1(n7399), .IN2(n7385), .IN3(n7513), .IN4(n7148), .Q(
        \U3/U92/Z_8 ) );
  AO22X1 U7574 ( .IN1(n7399), .IN2(n7148), .IN3(n7513), .IN4(n7314), .Q(
        \U3/U92/Z_7 ) );
  AO22X1 U7575 ( .IN1(n7399), .IN2(n7314), .IN3(n7513), .IN4(n7319), .Q(
        \U3/U92/Z_6 ) );
  AO22X1 U7576 ( .IN1(n7399), .IN2(n7319), .IN3(n7513), .IN4(n7324), .Q(
        \U3/U92/Z_5 ) );
  AO22X1 U7577 ( .IN1(n7399), .IN2(n7324), .IN3(n7513), .IN4(n7330), .Q(
        \U3/U92/Z_4 ) );
  AO22X1 U7578 ( .IN1(n7399), .IN2(n7330), .IN3(n7513), .IN4(n7332), .Q(
        \U3/U92/Z_3 ) );
  AO221X1 U7579 ( .IN1(n7513), .IN2(n7334), .IN3(n8000), .IN4(n7330), .IN5(
        n8001), .Q(\U3/U92/Z_2 ) );
  OAI21X1 U7580 ( .IN1(n7782), .IN2(n3714), .IN3(n8002), .QN(n8001) );
  INVX0 U7581 ( .INP(n7884), .ZN(n7513) );
  NOR2X0 U7582 ( .IN1(n3704), .IN2(n7782), .QN(\U3/U92/Z_11 ) );
  NOR2X0 U7583 ( .IN1(n3705), .IN2(n7782), .QN(\U3/U92/Z_10 ) );
  AO221X1 U7584 ( .IN1(n8003), .IN2(n7332), .IN3(n7399), .IN4(n7334), .IN5(
        n8004), .Q(\U3/U92/Z_1 ) );
  AO21X1 U7585 ( .IN1(n3723), .IN2(n3719), .IN3(n7799), .Q(n8003) );
  INVX0 U7586 ( .INP(n7869), .ZN(n7799) );
  AND2X1 U7587 ( .IN1(n7334), .IN2(n8000), .Q(\U3/U92/Z_0 ) );
  AO221X1 U7588 ( .IN1(n8005), .IN2(SP[9]), .IN3(n8004), .IN4(ID_PC[9]), .IN5(
        n8006), .Q(\U3/U91/Z_9 ) );
  AO22X1 U7589 ( .IN1(n9104), .IN2(n7399), .IN3(n8000), .IN4(n7173), .Q(n8006)
         );
  INVX0 U7590 ( .INP(n3684), .ZN(n7173) );
  AO221X1 U7591 ( .IN1(n8005), .IN2(SP[8]), .IN3(n8004), .IN4(ID_PC[8]), .IN5(
        n8007), .Q(\U3/U91/Z_8 ) );
  AO22X1 U7592 ( .IN1(n9106), .IN2(n7399), .IN3(n8000), .IN4(n7171), .Q(n8007)
         );
  INVX0 U7593 ( .INP(n3685), .ZN(n7171) );
  AO221X1 U7594 ( .IN1(n8005), .IN2(SP[7]), .IN3(n8004), .IN4(ID_PC[7]), .IN5(
        n8008), .Q(\U3/U91/Z_7 ) );
  AO22X1 U7595 ( .IN1(n9108), .IN2(n7399), .IN3(n8000), .IN4(n7169), .Q(n8008)
         );
  INVX0 U7596 ( .INP(n3686), .ZN(n7169) );
  AO221X1 U7597 ( .IN1(n8005), .IN2(SP[6]), .IN3(n8004), .IN4(ID_PC[6]), .IN5(
        n8009), .Q(\U3/U91/Z_6 ) );
  AO22X1 U7598 ( .IN1(n9110), .IN2(n7399), .IN3(n8000), .IN4(n7167), .Q(n8009)
         );
  INVX0 U7599 ( .INP(n3687), .ZN(n7167) );
  AO221X1 U7600 ( .IN1(n8005), .IN2(SP[5]), .IN3(n8004), .IN4(ID_PC[5]), .IN5(
        n8010), .Q(\U3/U91/Z_5 ) );
  AO22X1 U7601 ( .IN1(n9112), .IN2(n7399), .IN3(n8000), .IN4(n7165), .Q(n8010)
         );
  INVX0 U7602 ( .INP(n3688), .ZN(n7165) );
  AO221X1 U7603 ( .IN1(n8005), .IN2(SP[4]), .IN3(n8004), .IN4(ID_PC[4]), .IN5(
        n8011), .Q(\U3/U91/Z_4 ) );
  AO22X1 U7604 ( .IN1(n9114), .IN2(n7399), .IN3(n8000), .IN4(n7163), .Q(n8011)
         );
  INVX0 U7605 ( .INP(n3689), .ZN(n7163) );
  AO221X1 U7606 ( .IN1(n8005), .IN2(SP[31]), .IN3(n8004), .IN4(ID_PC[31]), 
        .IN5(n8012), .Q(\U3/U91/Z_31 ) );
  AO22X1 U7607 ( .IN1(n9028), .IN2(n7399), .IN3(n8000), .IN4(n7217), .Q(n8012)
         );
  INVX0 U7608 ( .INP(n3662), .ZN(n7217) );
  AO221X1 U7609 ( .IN1(n8005), .IN2(SP[30]), .IN3(n8004), .IN4(ID_PC[30]), 
        .IN5(n8013), .Q(\U3/U91/Z_30 ) );
  AO22X1 U7610 ( .IN1(n9062), .IN2(n7399), .IN3(n8000), .IN4(n7215), .Q(n8013)
         );
  INVX0 U7611 ( .INP(n3663), .ZN(n7215) );
  AO221X1 U7612 ( .IN1(n8005), .IN2(SP[3]), .IN3(n8004), .IN4(ID_PC[3]), .IN5(
        n8014), .Q(\U3/U91/Z_3 ) );
  AO22X1 U7613 ( .IN1(n9116), .IN2(n7399), .IN3(n8000), .IN4(n7161), .Q(n8014)
         );
  INVX0 U7614 ( .INP(n3690), .ZN(n7161) );
  AO221X1 U7615 ( .IN1(n8005), .IN2(SP[29]), .IN3(n8004), .IN4(ID_PC[29]), 
        .IN5(n8015), .Q(\U3/U91/Z_29 ) );
  AO22X1 U7616 ( .IN1(n9064), .IN2(n7399), .IN3(n8000), .IN4(n7213), .Q(n8015)
         );
  INVX0 U7617 ( .INP(n3664), .ZN(n7213) );
  AO221X1 U7618 ( .IN1(n8005), .IN2(SP[28]), .IN3(n8004), .IN4(ID_PC[28]), 
        .IN5(n8016), .Q(\U3/U91/Z_28 ) );
  AO22X1 U7619 ( .IN1(n9066), .IN2(n7399), .IN3(n8000), .IN4(n7211), .Q(n8016)
         );
  INVX0 U7620 ( .INP(n3665), .ZN(n7211) );
  AO221X1 U7621 ( .IN1(n8005), .IN2(SP[27]), .IN3(n8004), .IN4(ID_PC[27]), 
        .IN5(n8017), .Q(\U3/U91/Z_27 ) );
  AO22X1 U7622 ( .IN1(n9068), .IN2(n7399), .IN3(n8000), .IN4(n7209), .Q(n8017)
         );
  INVX0 U7623 ( .INP(n3666), .ZN(n7209) );
  AO221X1 U7624 ( .IN1(n8005), .IN2(SP[26]), .IN3(n8004), .IN4(ID_PC[26]), 
        .IN5(n8018), .Q(\U3/U91/Z_26 ) );
  AO22X1 U7625 ( .IN1(n9070), .IN2(n7399), .IN3(n8000), .IN4(n7207), .Q(n8018)
         );
  INVX0 U7626 ( .INP(n3667), .ZN(n7207) );
  AO221X1 U7627 ( .IN1(n8005), .IN2(SP[25]), .IN3(n8004), .IN4(ID_PC[25]), 
        .IN5(n8019), .Q(\U3/U91/Z_25 ) );
  AO22X1 U7628 ( .IN1(n9072), .IN2(n7399), .IN3(n8000), .IN4(n7205), .Q(n8019)
         );
  INVX0 U7629 ( .INP(n3668), .ZN(n7205) );
  AO221X1 U7630 ( .IN1(n8005), .IN2(SP[24]), .IN3(n8004), .IN4(ID_PC[24]), 
        .IN5(n8020), .Q(\U3/U91/Z_24 ) );
  AO22X1 U7631 ( .IN1(n9074), .IN2(n7399), .IN3(n8000), .IN4(n7203), .Q(n8020)
         );
  INVX0 U7632 ( .INP(n3669), .ZN(n7203) );
  AO221X1 U7633 ( .IN1(n8005), .IN2(SP[23]), .IN3(n8004), .IN4(ID_PC[23]), 
        .IN5(n8021), .Q(\U3/U91/Z_23 ) );
  AO22X1 U7634 ( .IN1(n9076), .IN2(n7399), .IN3(n8000), .IN4(n7201), .Q(n8021)
         );
  INVX0 U7635 ( .INP(n3670), .ZN(n7201) );
  AO221X1 U7636 ( .IN1(n8005), .IN2(SP[22]), .IN3(n8004), .IN4(ID_PC[22]), 
        .IN5(n8022), .Q(\U3/U91/Z_22 ) );
  AO22X1 U7637 ( .IN1(n9078), .IN2(n7399), .IN3(n8000), .IN4(n7199), .Q(n8022)
         );
  INVX0 U7638 ( .INP(n3671), .ZN(n7199) );
  AO221X1 U7639 ( .IN1(n8005), .IN2(SP[21]), .IN3(n8004), .IN4(ID_PC[21]), 
        .IN5(n8023), .Q(\U3/U91/Z_21 ) );
  AO22X1 U7640 ( .IN1(n9080), .IN2(n7399), .IN3(n8000), .IN4(n7197), .Q(n8023)
         );
  INVX0 U7641 ( .INP(n3672), .ZN(n7197) );
  AO221X1 U7642 ( .IN1(n8005), .IN2(SP[20]), .IN3(n8004), .IN4(ID_PC[20]), 
        .IN5(n8024), .Q(\U3/U91/Z_20 ) );
  AO22X1 U7643 ( .IN1(n9082), .IN2(n7399), .IN3(n8000), .IN4(n7195), .Q(n8024)
         );
  INVX0 U7644 ( .INP(n3673), .ZN(n7195) );
  AO221X1 U7645 ( .IN1(n8005), .IN2(SP[2]), .IN3(n8004), .IN4(ID_PC[2]), .IN5(
        n8025), .Q(\U3/U91/Z_2 ) );
  AO22X1 U7646 ( .IN1(n9118), .IN2(n7399), .IN3(n8000), .IN4(n7159), .Q(n8025)
         );
  INVX0 U7647 ( .INP(n3691), .ZN(n7159) );
  AO221X1 U7648 ( .IN1(n8005), .IN2(SP[19]), .IN3(n8004), .IN4(ID_PC[19]), 
        .IN5(n8026), .Q(\U3/U91/Z_19 ) );
  AO22X1 U7649 ( .IN1(n9084), .IN2(n7399), .IN3(n8000), .IN4(n7193), .Q(n8026)
         );
  INVX0 U7650 ( .INP(n3674), .ZN(n7193) );
  AO221X1 U7651 ( .IN1(n8005), .IN2(SP[18]), .IN3(n8004), .IN4(ID_PC[18]), 
        .IN5(n8027), .Q(\U3/U91/Z_18 ) );
  AO22X1 U7652 ( .IN1(n9086), .IN2(n7399), .IN3(n8000), .IN4(n7191), .Q(n8027)
         );
  INVX0 U7653 ( .INP(n3675), .ZN(n7191) );
  AO221X1 U7654 ( .IN1(n8005), .IN2(SP[17]), .IN3(n8004), .IN4(ID_PC[17]), 
        .IN5(n8028), .Q(\U3/U91/Z_17 ) );
  AO22X1 U7655 ( .IN1(n9088), .IN2(n7399), .IN3(n8000), .IN4(n7189), .Q(n8028)
         );
  INVX0 U7656 ( .INP(n3676), .ZN(n7189) );
  AO221X1 U7657 ( .IN1(n8005), .IN2(SP[16]), .IN3(n8004), .IN4(ID_PC[16]), 
        .IN5(n8029), .Q(\U3/U91/Z_16 ) );
  AO22X1 U7658 ( .IN1(n9090), .IN2(n7399), .IN3(n8000), .IN4(n7187), .Q(n8029)
         );
  INVX0 U7659 ( .INP(n3677), .ZN(n7187) );
  AO221X1 U7660 ( .IN1(n8005), .IN2(SP[15]), .IN3(n8004), .IN4(ID_PC[15]), 
        .IN5(n8030), .Q(\U3/U91/Z_15 ) );
  AO22X1 U7661 ( .IN1(n9092), .IN2(n7399), .IN3(n8000), .IN4(n7185), .Q(n8030)
         );
  INVX0 U7662 ( .INP(n3678), .ZN(n7185) );
  AO221X1 U7663 ( .IN1(n8005), .IN2(SP[14]), .IN3(n8004), .IN4(ID_PC[14]), 
        .IN5(n8031), .Q(\U3/U91/Z_14 ) );
  AO22X1 U7664 ( .IN1(n9094), .IN2(n7399), .IN3(n8000), .IN4(n7183), .Q(n8031)
         );
  INVX0 U7665 ( .INP(n3679), .ZN(n7183) );
  AO221X1 U7666 ( .IN1(n8005), .IN2(SP[13]), .IN3(n8004), .IN4(ID_PC[13]), 
        .IN5(n8032), .Q(\U3/U91/Z_13 ) );
  AO22X1 U7667 ( .IN1(n9096), .IN2(n7399), .IN3(n8000), .IN4(n7181), .Q(n8032)
         );
  INVX0 U7668 ( .INP(n3680), .ZN(n7181) );
  AO221X1 U7669 ( .IN1(n8005), .IN2(SP[12]), .IN3(n8004), .IN4(ID_PC[12]), 
        .IN5(n8033), .Q(\U3/U91/Z_12 ) );
  AO22X1 U7670 ( .IN1(n9098), .IN2(n7399), .IN3(n8000), .IN4(n7179), .Q(n8033)
         );
  INVX0 U7671 ( .INP(n3681), .ZN(n7179) );
  AO221X1 U7672 ( .IN1(n8005), .IN2(SP[11]), .IN3(n8004), .IN4(ID_PC[11]), 
        .IN5(n8034), .Q(\U3/U91/Z_11 ) );
  AO22X1 U7673 ( .IN1(n9100), .IN2(n7399), .IN3(n8000), .IN4(n7177), .Q(n8034)
         );
  INVX0 U7674 ( .INP(n3682), .ZN(n7177) );
  AO221X1 U7675 ( .IN1(n8005), .IN2(SP[10]), .IN3(n8004), .IN4(ID_PC[10]), 
        .IN5(n8035), .Q(\U3/U91/Z_10 ) );
  AO22X1 U7676 ( .IN1(n9102), .IN2(n7399), .IN3(n8000), .IN4(n7175), .Q(n8035)
         );
  INVX0 U7677 ( .INP(n3683), .ZN(n7175) );
  AO221X1 U7678 ( .IN1(n8005), .IN2(n7391), .IN3(n9171), .IN4(n8004), .IN5(
        n8036), .Q(\U3/U91/Z_1 ) );
  AO22X1 U7679 ( .IN1(n9120), .IN2(n7399), .IN3(n8000), .IN4(n7157), .Q(n8036)
         );
  INVX0 U7680 ( .INP(n3692), .ZN(n7157) );
  INVX0 U7681 ( .INP(n3573), .ZN(n7391) );
  AO221X1 U7682 ( .IN1(n8000), .IN2(n7155), .IN3(n7399), .IN4(n9170), .IN5(
        n8037), .Q(\U3/U91/Z_0 ) );
  AO22X1 U7683 ( .IN1(n9172), .IN2(n8004), .IN3(n8005), .IN4(n7390), .Q(n8037)
         );
  INVX0 U7684 ( .INP(n3574), .ZN(n7390) );
  NAND2X0 U7685 ( .IN1(n8002), .IN2(n7884), .QN(n8005) );
  NAND2X0 U7686 ( .IN1(\r1720/A[3] ), .IN2(n3723), .QN(n7884) );
  OA21X1 U7687 ( .IN1(n3721), .IN2(n3723), .IN3(n7579), .Q(n8002) );
  NAND2X0 U7688 ( .IN1(n7531), .IN2(n7800), .QN(n8004) );
  NAND2X0 U7689 ( .IN1(n7777), .IN2(n7512), .QN(n7800) );
  NAND2X0 U7690 ( .IN1(n3716), .IN2(n5695), .QN(n7531) );
  INVX0 U7691 ( .INP(n7782), .ZN(n7399) );
  INVX0 U7692 ( .INP(n3693), .ZN(n7155) );
  NAND2X0 U7693 ( .IN1(n7870), .IN2(n7869), .QN(n8000) );
  NOR2X0 U7694 ( .IN1(n7499), .IN2(n4486), .QN(\U3/U89/Z_0 ) );
  AO221X1 U7695 ( .IN1(n8038), .IN2(n7276), .IN3(n7777), .IN4(ID_imm_offset[8]), .IN5(n8039), .Q(\U3/U88/Z_9 ) );
  AO22X1 U7696 ( .IN1(n8040), .IN2(n7385), .IN3(n8038), .IN4(n7275), .Q(
        \U3/U88/Z_8 ) );
  AO222X1 U7697 ( .IN1(n7400), .IN2(n7385), .IN3(n8038), .IN4(n7274), .IN5(
        n8040), .IN6(n7148), .Q(\U3/U88/Z_7 ) );
  AO222X1 U7698 ( .IN1(n7400), .IN2(n7148), .IN3(n8038), .IN4(n7273), .IN5(
        n8040), .IN6(n7314), .Q(\U3/U88/Z_6 ) );
  AO222X1 U7699 ( .IN1(n7400), .IN2(n7314), .IN3(n8038), .IN4(n7272), .IN5(
        n8040), .IN6(n7319), .Q(\U3/U88/Z_5 ) );
  AO222X1 U7700 ( .IN1(n7400), .IN2(n7319), .IN3(n8038), .IN4(n7271), .IN5(
        n8040), .IN6(n7324), .Q(\U3/U88/Z_4 ) );
  NOR2X0 U7701 ( .IN1(n4454), .IN2(n7508), .QN(\U3/U88/Z_32 ) );
  AO21X1 U7702 ( .IN1(n8038), .IN2(n7298), .IN3(n8041), .Q(\U3/U88/Z_31 ) );
  AO21X1 U7703 ( .IN1(n8038), .IN2(n7297), .IN3(n8041), .Q(\U3/U88/Z_30 ) );
  AO222X1 U7704 ( .IN1(n7400), .IN2(n7324), .IN3(n8038), .IN4(n7270), .IN5(
        n8040), .IN6(n7330), .Q(\U3/U88/Z_3 ) );
  AO21X1 U7705 ( .IN1(n8038), .IN2(n7296), .IN3(n8041), .Q(\U3/U88/Z_29 ) );
  AO21X1 U7706 ( .IN1(n8038), .IN2(n7295), .IN3(n8041), .Q(\U3/U88/Z_28 ) );
  AO21X1 U7707 ( .IN1(n8038), .IN2(n7294), .IN3(n8041), .Q(\U3/U88/Z_27 ) );
  AO21X1 U7708 ( .IN1(n8038), .IN2(n7293), .IN3(n8041), .Q(\U3/U88/Z_26 ) );
  AO21X1 U7709 ( .IN1(n8038), .IN2(n7292), .IN3(n8041), .Q(\U3/U88/Z_25 ) );
  AO21X1 U7710 ( .IN1(n8038), .IN2(n7291), .IN3(n8041), .Q(\U3/U88/Z_24 ) );
  AO21X1 U7711 ( .IN1(n8038), .IN2(n7290), .IN3(n8041), .Q(\U3/U88/Z_23 ) );
  AO21X1 U7712 ( .IN1(n8038), .IN2(n7289), .IN3(n8041), .Q(\U3/U88/Z_22 ) );
  AO21X1 U7713 ( .IN1(n7770), .IN2(n7116), .IN3(n8042), .Q(n8041) );
  AO221X1 U7714 ( .IN1(n8038), .IN2(n7288), .IN3(n7770), .IN4(ID_imm_offset[9]), .IN5(n8042), .Q(\U3/U88/Z_21 ) );
  AO221X1 U7715 ( .IN1(n8038), .IN2(n7287), .IN3(n7770), .IN4(ID_imm_offset[8]), .IN5(n8042), .Q(\U3/U88/Z_20 ) );
  AO222X1 U7716 ( .IN1(n7400), .IN2(n7330), .IN3(n8038), .IN4(n7269), .IN5(
        n8040), .IN6(n7332), .Q(\U3/U88/Z_2 ) );
  AO221X1 U7717 ( .IN1(n8038), .IN2(n7286), .IN3(n7770), .IN4(n7385), .IN5(
        n8042), .Q(\U3/U88/Z_19 ) );
  INVX0 U7718 ( .INP(n3696), .ZN(n7385) );
  AO221X1 U7719 ( .IN1(n8038), .IN2(n7285), .IN3(n7770), .IN4(n7148), .IN5(
        n8042), .Q(\U3/U88/Z_18 ) );
  AO221X1 U7720 ( .IN1(n8038), .IN2(n7284), .IN3(n7770), .IN4(n7314), .IN5(
        n8042), .Q(\U3/U88/Z_17 ) );
  INVX0 U7721 ( .INP(n3629), .ZN(n7314) );
  AO221X1 U7722 ( .IN1(n8038), .IN2(n7283), .IN3(n7770), .IN4(n7319), .IN5(
        n8042), .Q(\U3/U88/Z_16 ) );
  AO221X1 U7723 ( .IN1(n8038), .IN2(n7282), .IN3(n7770), .IN4(n7324), .IN5(
        n8042), .Q(\U3/U88/Z_15 ) );
  INVX0 U7724 ( .INP(n3627), .ZN(n7324) );
  AO221X1 U7725 ( .IN1(n8038), .IN2(n7281), .IN3(n7770), .IN4(n7330), .IN5(
        n8042), .Q(\U3/U88/Z_14 ) );
  AO221X1 U7726 ( .IN1(n8038), .IN2(n7280), .IN3(n7770), .IN4(n7332), .IN5(
        n8042), .Q(\U3/U88/Z_13 ) );
  AO221X1 U7727 ( .IN1(n8038), .IN2(n7279), .IN3(n7770), .IN4(n7334), .IN5(
        n8042), .Q(\U3/U88/Z_12 ) );
  AO21X1 U7728 ( .IN1(n8038), .IN2(n7278), .IN3(n8042), .Q(\U3/U88/Z_11 ) );
  AO21X1 U7729 ( .IN1(n7777), .IN2(n7116), .IN3(n8039), .Q(n8042) );
  INVX0 U7730 ( .INP(n3704), .ZN(n7116) );
  AO221X1 U7731 ( .IN1(n8038), .IN2(n7277), .IN3(n7777), .IN4(ID_imm_offset[9]), .IN5(n8039), .Q(\U3/U88/Z_10 ) );
  NOR2X0 U7732 ( .IN1(n7458), .IN2(n3696), .QN(n8039) );
  INVX0 U7733 ( .INP(n7394), .ZN(n7777) );
  AO222X1 U7734 ( .IN1(n7400), .IN2(n7332), .IN3(n8038), .IN4(n7268), .IN5(
        n8040), .IN6(n7334), .Q(\U3/U88/Z_1 ) );
  INVX0 U7735 ( .INP(n3714), .ZN(n7332) );
  AO22X1 U7736 ( .IN1(n7400), .IN2(n7334), .IN3(n8038), .IN4(n7265), .Q(
        \U3/U88/Z_0 ) );
  OR2X1 U7737 ( .IN1(n7555), .IN2(\U3/U90/Z_0 ), .Q(n8038) );
  INVX0 U7738 ( .INP(n7499), .ZN(n7555) );
  INVX0 U7739 ( .INP(n3713), .ZN(n7334) );
  INVX0 U7740 ( .INP(n7556), .ZN(n7400) );
  AO222X1 U7741 ( .IN1(n8043), .IN2(n7254), .IN3(n7770), .IN4(ID_PC[9]), .IN5(
        n529), .IN6(n8040), .Q(\U3/U87/Z_9 ) );
  AO222X1 U7742 ( .IN1(n8043), .IN2(n7255), .IN3(n7770), .IN4(ID_PC[8]), .IN5(
        n530), .IN6(n8040), .Q(\U3/U87/Z_8 ) );
  AO222X1 U7743 ( .IN1(n8043), .IN2(n7256), .IN3(n7770), .IN4(ID_PC[7]), .IN5(
        n531), .IN6(n8040), .Q(\U3/U87/Z_7 ) );
  AO222X1 U7744 ( .IN1(n8043), .IN2(n7257), .IN3(n7770), .IN4(ID_PC[6]), .IN5(
        n532), .IN6(n8040), .Q(\U3/U87/Z_6 ) );
  AO222X1 U7745 ( .IN1(n8043), .IN2(n7258), .IN3(n7770), .IN4(ID_PC[5]), .IN5(
        n533), .IN6(n8040), .Q(\U3/U87/Z_5 ) );
  AO222X1 U7746 ( .IN1(n8043), .IN2(n7259), .IN3(n7770), .IN4(ID_PC[4]), .IN5(
        n534), .IN6(n8040), .Q(\U3/U87/Z_4 ) );
  AO222X1 U7747 ( .IN1(n8043), .IN2(n7232), .IN3(n7770), .IN4(ID_PC[31]), 
        .IN5(n507), .IN6(n8040), .Q(\U3/U87/Z_31 ) );
  AO222X1 U7748 ( .IN1(n8043), .IN2(n7233), .IN3(n7770), .IN4(ID_PC[30]), 
        .IN5(n508), .IN6(n8040), .Q(\U3/U87/Z_30 ) );
  AO222X1 U7749 ( .IN1(n8043), .IN2(n7260), .IN3(n7770), .IN4(ID_PC[3]), .IN5(
        n535), .IN6(n8040), .Q(\U3/U87/Z_3 ) );
  AO222X1 U7750 ( .IN1(n8043), .IN2(n7234), .IN3(n7770), .IN4(ID_PC[29]), 
        .IN5(n509), .IN6(n8040), .Q(\U3/U87/Z_29 ) );
  AO222X1 U7751 ( .IN1(n8043), .IN2(n7235), .IN3(n7770), .IN4(ID_PC[28]), 
        .IN5(n510), .IN6(n8040), .Q(\U3/U87/Z_28 ) );
  AO222X1 U7752 ( .IN1(n8043), .IN2(n7236), .IN3(n7770), .IN4(ID_PC[27]), 
        .IN5(n511), .IN6(n8040), .Q(\U3/U87/Z_27 ) );
  AO222X1 U7753 ( .IN1(n8043), .IN2(n7237), .IN3(n7770), .IN4(ID_PC[26]), 
        .IN5(n512), .IN6(n8040), .Q(\U3/U87/Z_26 ) );
  AO222X1 U7754 ( .IN1(n8043), .IN2(n7238), .IN3(n7770), .IN4(ID_PC[25]), 
        .IN5(n513), .IN6(n8040), .Q(\U3/U87/Z_25 ) );
  AO222X1 U7755 ( .IN1(n8043), .IN2(n7239), .IN3(n7770), .IN4(ID_PC[24]), 
        .IN5(n514), .IN6(n8040), .Q(\U3/U87/Z_24 ) );
  AO222X1 U7756 ( .IN1(n8043), .IN2(n7240), .IN3(n7770), .IN4(ID_PC[23]), 
        .IN5(n515), .IN6(n8040), .Q(\U3/U87/Z_23 ) );
  AO222X1 U7757 ( .IN1(n8043), .IN2(n7241), .IN3(n7770), .IN4(ID_PC[22]), 
        .IN5(n516), .IN6(n8040), .Q(\U3/U87/Z_22 ) );
  AO222X1 U7758 ( .IN1(n8043), .IN2(n7242), .IN3(n7770), .IN4(ID_PC[21]), 
        .IN5(n517), .IN6(n8040), .Q(\U3/U87/Z_21 ) );
  AO222X1 U7759 ( .IN1(n8043), .IN2(n7243), .IN3(n7770), .IN4(ID_PC[20]), 
        .IN5(n518), .IN6(n8040), .Q(\U3/U87/Z_20 ) );
  AO222X1 U7760 ( .IN1(n8043), .IN2(n7261), .IN3(n7770), .IN4(ID_PC[2]), .IN5(
        n536), .IN6(n8040), .Q(\U3/U87/Z_2 ) );
  AO222X1 U7761 ( .IN1(n8043), .IN2(n7244), .IN3(n7770), .IN4(ID_PC[19]), 
        .IN5(n519), .IN6(n8040), .Q(\U3/U87/Z_19 ) );
  AO222X1 U7762 ( .IN1(n8043), .IN2(n7245), .IN3(n7770), .IN4(ID_PC[18]), 
        .IN5(n520), .IN6(n8040), .Q(\U3/U87/Z_18 ) );
  AO222X1 U7763 ( .IN1(n8043), .IN2(n7246), .IN3(n7770), .IN4(ID_PC[17]), 
        .IN5(n521), .IN6(n8040), .Q(\U3/U87/Z_17 ) );
  AO222X1 U7764 ( .IN1(n8043), .IN2(n7247), .IN3(n7770), .IN4(ID_PC[16]), 
        .IN5(n522), .IN6(n8040), .Q(\U3/U87/Z_16 ) );
  AO222X1 U7765 ( .IN1(n8043), .IN2(n7248), .IN3(n7770), .IN4(ID_PC[15]), 
        .IN5(n523), .IN6(n8040), .Q(\U3/U87/Z_15 ) );
  AO222X1 U7766 ( .IN1(n8043), .IN2(n7249), .IN3(n7770), .IN4(ID_PC[14]), 
        .IN5(n524), .IN6(n8040), .Q(\U3/U87/Z_14 ) );
  AO222X1 U7767 ( .IN1(n8043), .IN2(n7250), .IN3(n7770), .IN4(ID_PC[13]), 
        .IN5(n525), .IN6(n8040), .Q(\U3/U87/Z_13 ) );
  AO222X1 U7768 ( .IN1(n8043), .IN2(n7251), .IN3(n7770), .IN4(ID_PC[12]), 
        .IN5(n526), .IN6(n8040), .Q(\U3/U87/Z_12 ) );
  AO222X1 U7769 ( .IN1(n8043), .IN2(n7252), .IN3(n7770), .IN4(ID_PC[11]), 
        .IN5(n527), .IN6(n8040), .Q(\U3/U87/Z_11 ) );
  AO222X1 U7770 ( .IN1(n8043), .IN2(n7253), .IN3(n7770), .IN4(ID_PC[10]), 
        .IN5(n528), .IN6(n8040), .Q(\U3/U87/Z_10 ) );
  AO222X1 U7771 ( .IN1(n8043), .IN2(n7262), .IN3(n9171), .IN4(n7770), .IN5(
        n537), .IN6(n8040), .Q(\U3/U87/Z_1 ) );
  AO222X1 U7772 ( .IN1(n8043), .IN2(n7263), .IN3(n9172), .IN4(n7770), .IN5(
        n538), .IN6(n8040), .Q(\U3/U87/Z_0 ) );
  NAND2X0 U7773 ( .IN1(n7394), .IN2(n7458), .QN(n8040) );
  NAND3X0 U7774 ( .IN1(\r1720/A[3] ), .IN2(n7521), .IN3(n3716), .QN(n7458) );
  INVX0 U7775 ( .INP(n7797), .ZN(n7770) );
  NAND2X0 U7776 ( .IN1(n7784), .IN2(n7521), .QN(n7797) );
  INVX0 U7777 ( .INP(n7395), .ZN(n7784) );
  NAND2X0 U7778 ( .IN1(n7526), .IN2(n7447), .QN(n7395) );
  NAND3X0 U7779 ( .IN1(n7556), .IN2(n7782), .IN3(n7499), .QN(n8043) );
  NAND2X0 U7780 ( .IN1(n3716), .IN2(n3723), .QN(n7499) );
  NAND2X0 U7781 ( .IN1(\r1720/A[3] ), .IN2(n7447), .QN(n7782) );
  NAND2X0 U7782 ( .IN1(n3719), .IN2(n5695), .QN(n7556) );
  AO21X1 U7783 ( .IN1(n8044), .IN2(n7384), .IN3(n9191), .Q(N6325) );
  NAND2X0 U7784 ( .IN1(n8045), .IN2(n7889), .QN(n7384) );
  OA222X1 U7785 ( .IN1(n7869), .IN2(\r1720/A[3] ), .IN3(n8046), .IN4(n3719), 
        .IN5(n7508), .IN6(n3723), .Q(n7889) );
  NAND2X0 U7786 ( .IN1(n3723), .IN2(n7447), .QN(n7869) );
  MUX21X1 U7787 ( .IN1(n7450), .IN2(n7545), .S(n3719), .Q(n8045) );
  INVX0 U7788 ( .INP(n7457), .ZN(n7545) );
  NAND2X0 U7789 ( .IN1(n5696), .IN2(n7512), .QN(n7457) );
  INVX0 U7790 ( .INP(n3720), .ZN(n7512) );
  OR3X1 U7791 ( .IN1(n7394), .IN2(n3721), .IN3(n7579), .Q(n8044) );
  NAND3X0 U7792 ( .IN1(n3720), .IN2(n7521), .IN3(n3723), .QN(n7579) );
  NAND2X0 U7793 ( .IN1(n3716), .IN2(n7526), .QN(n7394) );
  AO21X1 U7794 ( .IN1(n8047), .IN2(n8048), .IN3(n9191), .Q(N6323) );
  NAND3X0 U7795 ( .IN1(n7549), .IN2(n7870), .IN3(n7576), .QN(n8048) );
  NOR2X0 U7796 ( .IN1(n5753), .IN2(n3720), .QN(n7576) );
  NAND2X0 U7797 ( .IN1(n3716), .IN2(n3719), .QN(n7870) );
  NAND2X0 U7798 ( .IN1(n8046), .IN2(n7521), .QN(n7549) );
  INVX0 U7799 ( .INP(n3719), .ZN(n7521) );
  NOR2X0 U7800 ( .IN1(n3723), .IN2(n3716), .QN(n8046) );
  NAND3X0 U7801 ( .IN1(n7501), .IN2(n7450), .IN3(n7451), .QN(n8047) );
  INVX0 U7802 ( .INP(n7806), .ZN(n7451) );
  NAND2X0 U7803 ( .IN1(n7526), .IN2(n5695), .QN(n7806) );
  INVX0 U7804 ( .INP(n7550), .ZN(n7450) );
  NAND2X0 U7805 ( .IN1(n3720), .IN2(n5696), .QN(n7550) );
  INVX0 U7806 ( .INP(n7508), .ZN(n7501) );
  NAND2X0 U7807 ( .IN1(n3719), .IN2(n7447), .QN(n7508) );
  INVX0 U7808 ( .INP(n3716), .ZN(n7447) );
  NAND2X0 U7809 ( .IN1(n3630), .IN2(n4485), .QN(N5077) );
  NAND2X0 U7810 ( .IN1(n3631), .IN2(n4484), .QN(N5076) );
  NAND2X0 U7811 ( .IN1(n3632), .IN2(n4483), .QN(N5075) );
  NAND2X0 U7812 ( .IN1(n3633), .IN2(n4482), .QN(N5074) );
  NAND2X0 U7813 ( .IN1(n3634), .IN2(n4481), .QN(N5073) );
  NAND2X0 U7814 ( .IN1(n3635), .IN2(n4480), .QN(N5072) );
  NAND2X0 U7815 ( .IN1(n3636), .IN2(n4479), .QN(N5071) );
  NAND2X0 U7816 ( .IN1(n3637), .IN2(n4478), .QN(N5070) );
  NAND2X0 U7817 ( .IN1(n4477), .IN2(n3638), .QN(N5069) );
  NAND2X0 U7818 ( .IN1(n4476), .IN2(n3639), .QN(N5068) );
  NAND2X0 U7819 ( .IN1(n4475), .IN2(n3640), .QN(N5067) );
  NAND2X0 U7820 ( .IN1(n4474), .IN2(n3641), .QN(N5066) );
  NAND2X0 U7821 ( .IN1(n4473), .IN2(n3642), .QN(N5065) );
  NAND2X0 U7822 ( .IN1(n4472), .IN2(n3643), .QN(N5064) );
  NAND2X0 U7823 ( .IN1(n4471), .IN2(n3644), .QN(N5063) );
  NAND2X0 U7824 ( .IN1(n4470), .IN2(n3645), .QN(N5062) );
  NAND2X0 U7825 ( .IN1(n4469), .IN2(n3646), .QN(N5061) );
  NAND2X0 U7826 ( .IN1(n4468), .IN2(n3647), .QN(N5060) );
  NAND2X0 U7827 ( .IN1(n4467), .IN2(n3648), .QN(N5059) );
  NAND2X0 U7828 ( .IN1(n4466), .IN2(n3649), .QN(N5058) );
  NAND2X0 U7829 ( .IN1(n4465), .IN2(n3650), .QN(N5057) );
  NAND2X0 U7830 ( .IN1(n4464), .IN2(n3651), .QN(N5056) );
  NAND2X0 U7831 ( .IN1(n4463), .IN2(n3652), .QN(N5055) );
  NAND2X0 U7832 ( .IN1(n4462), .IN2(n3653), .QN(N5054) );
  NAND2X0 U7833 ( .IN1(n4461), .IN2(n3654), .QN(N5053) );
  NAND2X0 U7834 ( .IN1(n4460), .IN2(n3655), .QN(N5052) );
  NAND2X0 U7835 ( .IN1(n4459), .IN2(n3656), .QN(N5051) );
  NAND2X0 U7836 ( .IN1(n4458), .IN2(n3657), .QN(N5050) );
  NAND2X0 U7837 ( .IN1(n4457), .IN2(n3658), .QN(N5049) );
  NAND2X0 U7838 ( .IN1(n4456), .IN2(n3659), .QN(N5048) );
  NAND2X0 U7839 ( .IN1(n4455), .IN2(n3660), .QN(N5047) );
  NAND2X0 U7840 ( .IN1(n4454), .IN2(n3661), .QN(N5046) );
  AND2X1 U7841 ( .IN1(N4947), .IN2(n7769), .Q(N4979) );
  AND2X1 U7842 ( .IN1(N4946), .IN2(n7769), .Q(N4978) );
  AND2X1 U7843 ( .IN1(N4945), .IN2(n7769), .Q(N4977) );
  AND2X1 U7844 ( .IN1(N4944), .IN2(n7769), .Q(N4976) );
  AND2X1 U7845 ( .IN1(N4943), .IN2(n7769), .Q(N4975) );
  AND2X1 U7846 ( .IN1(N4942), .IN2(n7769), .Q(N4974) );
  AND2X1 U7847 ( .IN1(N4941), .IN2(n7769), .Q(N4973) );
  AND2X1 U7848 ( .IN1(N4940), .IN2(n7769), .Q(N4972) );
  AND2X1 U7849 ( .IN1(N4939), .IN2(n7769), .Q(N4971) );
  AND2X1 U7850 ( .IN1(N4938), .IN2(n7769), .Q(N4970) );
  AND2X1 U7851 ( .IN1(N4937), .IN2(n7769), .Q(N4969) );
  AND2X1 U7852 ( .IN1(N4936), .IN2(n7769), .Q(N4968) );
  AND2X1 U7853 ( .IN1(N4935), .IN2(n7769), .Q(N4967) );
  AND2X1 U7854 ( .IN1(N4934), .IN2(n7769), .Q(N4966) );
  AND2X1 U7855 ( .IN1(N4933), .IN2(n7769), .Q(N4965) );
  AND2X1 U7856 ( .IN1(N4932), .IN2(n7769), .Q(N4964) );
  AND2X1 U7857 ( .IN1(N4931), .IN2(n7769), .Q(N4963) );
  AND2X1 U7858 ( .IN1(N4930), .IN2(n7769), .Q(N4962) );
  AND2X1 U7859 ( .IN1(N4929), .IN2(n7769), .Q(N4961) );
  AND2X1 U7860 ( .IN1(N4928), .IN2(n7769), .Q(N4960) );
  AND2X1 U7861 ( .IN1(N4927), .IN2(n7769), .Q(N4959) );
  AND2X1 U7862 ( .IN1(N4926), .IN2(n7769), .Q(N4958) );
  AND2X1 U7863 ( .IN1(N4925), .IN2(n7769), .Q(N4957) );
  AND2X1 U7864 ( .IN1(N4924), .IN2(n7769), .Q(N4956) );
  AND2X1 U7865 ( .IN1(N4923), .IN2(n7769), .Q(N4955) );
  AND2X1 U7866 ( .IN1(N4922), .IN2(n7769), .Q(N4954) );
  AND2X1 U7867 ( .IN1(N4921), .IN2(n7769), .Q(N4953) );
  AND2X1 U7868 ( .IN1(N4920), .IN2(n7769), .Q(N4952) );
  AND2X1 U7869 ( .IN1(N4919), .IN2(n7769), .Q(N4951) );
  AND2X1 U7870 ( .IN1(N4918), .IN2(n7769), .Q(N4950) );
  AND2X1 U7871 ( .IN1(N4917), .IN2(n7769), .Q(N4949) );
  AND2X1 U7872 ( .IN1(N4916), .IN2(n7769), .Q(N4948) );
  AND2X1 U7873 ( .IN1(N4844), .IN2(n7769), .Q(N4877) );
  AND2X1 U7874 ( .IN1(N4843), .IN2(n7769), .Q(N4876) );
  AND2X1 U7875 ( .IN1(N4842), .IN2(n7769), .Q(N4875) );
  AND2X1 U7876 ( .IN1(N4841), .IN2(n7769), .Q(N4874) );
  AND2X1 U7877 ( .IN1(N4840), .IN2(n7769), .Q(N4873) );
  AND2X1 U7878 ( .IN1(N4839), .IN2(n7769), .Q(N4872) );
  AND2X1 U7879 ( .IN1(N4838), .IN2(n7769), .Q(N4871) );
  AND2X1 U7880 ( .IN1(N4837), .IN2(n7769), .Q(N4870) );
  AND2X1 U7881 ( .IN1(N4836), .IN2(n7769), .Q(N4869) );
  AND2X1 U7882 ( .IN1(N4835), .IN2(n7769), .Q(N4868) );
  AND2X1 U7883 ( .IN1(N4834), .IN2(n7769), .Q(N4867) );
  AND2X1 U7884 ( .IN1(N4833), .IN2(n7769), .Q(N4866) );
  AND2X1 U7885 ( .IN1(N4832), .IN2(n7769), .Q(N4865) );
  AND2X1 U7886 ( .IN1(N4831), .IN2(n7769), .Q(N4864) );
  AND2X1 U7887 ( .IN1(N4830), .IN2(n7769), .Q(N4863) );
  AND2X1 U7888 ( .IN1(N4829), .IN2(n7769), .Q(N4862) );
  AND2X1 U7889 ( .IN1(N4828), .IN2(n7769), .Q(N4861) );
  AND2X1 U7890 ( .IN1(N4827), .IN2(n7769), .Q(N4860) );
  AND2X1 U7891 ( .IN1(N4826), .IN2(n7769), .Q(N4859) );
  AND2X1 U7892 ( .IN1(N4825), .IN2(n7769), .Q(N4858) );
  AND2X1 U7893 ( .IN1(N4824), .IN2(n7769), .Q(N4857) );
  AND2X1 U7894 ( .IN1(N4823), .IN2(n7769), .Q(N4856) );
  AND2X1 U7895 ( .IN1(N4822), .IN2(n7769), .Q(N4855) );
  AND2X1 U7896 ( .IN1(N4821), .IN2(n7769), .Q(N4854) );
  AND2X1 U7897 ( .IN1(N4820), .IN2(n7769), .Q(N4853) );
  AND2X1 U7898 ( .IN1(N4819), .IN2(n7769), .Q(N4852) );
  AND2X1 U7899 ( .IN1(N4818), .IN2(n7769), .Q(N4851) );
  AND2X1 U7900 ( .IN1(N4817), .IN2(n7769), .Q(N4850) );
  AND2X1 U7901 ( .IN1(N4816), .IN2(n7769), .Q(N4849) );
  AND2X1 U7902 ( .IN1(N4815), .IN2(n7769), .Q(N4848) );
  AND2X1 U7903 ( .IN1(N4814), .IN2(n7769), .Q(N4847) );
  AND2X1 U7904 ( .IN1(N4813), .IN2(n7769), .Q(N4846) );
  AOI22X1 U7905 ( .IN1(n7272), .IN2(n7875), .IN3(n8049), .IN4(n8050), .QN(
        n7769) );
  NAND3X0 U7906 ( .IN1(n4479), .IN2(n4478), .IN3(n4481), .QN(n8050) );
  NAND4X0 U7907 ( .IN1(n4485), .IN2(n4484), .IN3(n4483), .IN4(n4482), .QN(
        n7875) );
  MUX21X1 U7908 ( .IN1(N354), .IN2(n9061), .S(n9191), .Q(N466) );
  MUX21X1 U7909 ( .IN1(N353), .IN2(n9063), .S(n9191), .Q(N465) );
  MUX21X1 U7910 ( .IN1(N352), .IN2(n9065), .S(n9191), .Q(N464) );
  MUX21X1 U7911 ( .IN1(N351), .IN2(n9067), .S(n9191), .Q(N463) );
  MUX21X1 U7912 ( .IN1(N350), .IN2(n9069), .S(n9191), .Q(N462) );
  MUX21X1 U7913 ( .IN1(N349), .IN2(n9071), .S(n9191), .Q(N461) );
  MUX21X1 U7914 ( .IN1(N348), .IN2(n9073), .S(n9191), .Q(N460) );
  MUX21X1 U7915 ( .IN1(N347), .IN2(n9075), .S(n9191), .Q(N459) );
  MUX21X1 U7916 ( .IN1(N346), .IN2(n9077), .S(n9191), .Q(N458) );
  AO21X1 U7917 ( .IN1(n3630), .IN2(n7265), .IN3(N4382), .Q(N4578) );
  AO21X1 U7918 ( .IN1(n3631), .IN2(n7268), .IN3(N4381), .Q(N4577) );
  AO21X1 U7919 ( .IN1(n3632), .IN2(n7269), .IN3(N4380), .Q(N4576) );
  AO21X1 U7920 ( .IN1(n3633), .IN2(n7270), .IN3(N4379), .Q(N4575) );
  AO21X1 U7921 ( .IN1(n3634), .IN2(n7271), .IN3(N4378), .Q(N4574) );
  AO21X1 U7922 ( .IN1(n3635), .IN2(n7272), .IN3(N4377), .Q(N4573) );
  AO21X1 U7923 ( .IN1(n3636), .IN2(n7273), .IN3(N4376), .Q(N4572) );
  AO21X1 U7924 ( .IN1(n3637), .IN2(n7274), .IN3(N4375), .Q(N4571) );
  AO21X1 U7925 ( .IN1(n3638), .IN2(n7275), .IN3(N4374), .Q(N4570) );
  MUX21X1 U7926 ( .IN1(N345), .IN2(n9079), .S(n9191), .Q(N457) );
  AO21X1 U7927 ( .IN1(n3639), .IN2(n7276), .IN3(N4373), .Q(N4569) );
  AO21X1 U7928 ( .IN1(n3640), .IN2(n7277), .IN3(N4372), .Q(N4568) );
  AO21X1 U7929 ( .IN1(n3641), .IN2(n7278), .IN3(N4371), .Q(N4567) );
  AO21X1 U7930 ( .IN1(n3642), .IN2(n7279), .IN3(N4370), .Q(N4566) );
  AO21X1 U7931 ( .IN1(n3643), .IN2(n7280), .IN3(N4369), .Q(N4565) );
  AO21X1 U7932 ( .IN1(n3644), .IN2(n7281), .IN3(N4368), .Q(N4564) );
  AO21X1 U7933 ( .IN1(n3645), .IN2(n7282), .IN3(N4367), .Q(N4563) );
  AO21X1 U7934 ( .IN1(n3646), .IN2(n7283), .IN3(N4366), .Q(N4562) );
  AO21X1 U7935 ( .IN1(n3647), .IN2(n7284), .IN3(N4365), .Q(N4561) );
  AO21X1 U7936 ( .IN1(n3648), .IN2(n7285), .IN3(N4364), .Q(N4560) );
  MUX21X1 U7937 ( .IN1(N344), .IN2(n9081), .S(n9191), .Q(N456) );
  AO21X1 U7938 ( .IN1(n3649), .IN2(n7286), .IN3(N4363), .Q(N4559) );
  AO21X1 U7939 ( .IN1(n3650), .IN2(n7287), .IN3(N4362), .Q(N4558) );
  AO21X1 U7940 ( .IN1(n3651), .IN2(n7288), .IN3(N4361), .Q(N4557) );
  AO21X1 U7941 ( .IN1(n3652), .IN2(n7289), .IN3(N4360), .Q(N4556) );
  AO21X1 U7942 ( .IN1(n3653), .IN2(n7290), .IN3(N4359), .Q(N4555) );
  AO21X1 U7943 ( .IN1(n3654), .IN2(n7291), .IN3(N4358), .Q(N4554) );
  AO21X1 U7944 ( .IN1(n3655), .IN2(n7292), .IN3(N4357), .Q(N4553) );
  AO21X1 U7945 ( .IN1(n3656), .IN2(n7293), .IN3(N4356), .Q(N4552) );
  AO21X1 U7946 ( .IN1(n3657), .IN2(n7294), .IN3(N4355), .Q(N4551) );
  AO21X1 U7947 ( .IN1(n3658), .IN2(n7295), .IN3(N4354), .Q(N4550) );
  MUX21X1 U7948 ( .IN1(N343), .IN2(n9083), .S(n9191), .Q(N455) );
  AO21X1 U7949 ( .IN1(n3659), .IN2(n7296), .IN3(N4353), .Q(N4549) );
  AO21X1 U7950 ( .IN1(n3660), .IN2(n7297), .IN3(N4352), .Q(N4548) );
  AO21X1 U7951 ( .IN1(n3661), .IN2(n7298), .IN3(N4351), .Q(N4547) );
  MUX21X1 U7952 ( .IN1(N342), .IN2(n9085), .S(n9191), .Q(N454) );
  MUX21X1 U7953 ( .IN1(N341), .IN2(n9087), .S(n9191), .Q(N453) );
  MUX21X1 U7954 ( .IN1(N340), .IN2(n9089), .S(n9191), .Q(N452) );
  MUX21X1 U7955 ( .IN1(N339), .IN2(n9091), .S(n9191), .Q(N451) );
  MUX21X1 U7956 ( .IN1(N338), .IN2(n9093), .S(n9191), .Q(N450) );
  MUX21X1 U7957 ( .IN1(N337), .IN2(n9095), .S(n9191), .Q(N449) );
  MUX21X1 U7958 ( .IN1(N336), .IN2(n9097), .S(n9191), .Q(N448) );
  MUX21X1 U7959 ( .IN1(N335), .IN2(n9099), .S(n9191), .Q(N447) );
  MUX21X1 U7960 ( .IN1(N334), .IN2(n9101), .S(n9191), .Q(N446) );
  MUX21X1 U7961 ( .IN1(N333), .IN2(n9103), .S(n9191), .Q(N445) );
  MUX21X1 U7962 ( .IN1(N332), .IN2(n9105), .S(n9191), .Q(N444) );
  MUX21X1 U7963 ( .IN1(N331), .IN2(n9107), .S(n9191), .Q(N443) );
  MUX21X1 U7964 ( .IN1(N330), .IN2(n9109), .S(n9191), .Q(N442) );
  MUX21X1 U7965 ( .IN1(N329), .IN2(n9111), .S(n9191), .Q(N441) );
  MUX21X1 U7966 ( .IN1(N328), .IN2(n9113), .S(n9191), .Q(N440) );
  MUX21X1 U7967 ( .IN1(N327), .IN2(n9115), .S(n9191), .Q(N439) );
  NOR2X0 U7968 ( .IN1(n7265), .IN2(n3630), .QN(N4382) );
  INVX0 U7969 ( .INP(n4485), .ZN(n7265) );
  NOR2X0 U7970 ( .IN1(n7268), .IN2(n3631), .QN(N4381) );
  INVX0 U7971 ( .INP(n4484), .ZN(n7268) );
  NOR2X0 U7972 ( .IN1(n7269), .IN2(n3632), .QN(N4380) );
  INVX0 U7973 ( .INP(n4483), .ZN(n7269) );
  MUX21X1 U7974 ( .IN1(N326), .IN2(n9117), .S(n9191), .Q(N438) );
  NOR2X0 U7975 ( .IN1(n7270), .IN2(n3633), .QN(N4379) );
  INVX0 U7976 ( .INP(n4482), .ZN(n7270) );
  NOR2X0 U7977 ( .IN1(n7271), .IN2(n3634), .QN(N4378) );
  INVX0 U7978 ( .INP(n4481), .ZN(n7271) );
  NOR2X0 U7979 ( .IN1(n7272), .IN2(n3635), .QN(N4377) );
  INVX0 U7980 ( .INP(n4480), .ZN(n7272) );
  NOR2X0 U7981 ( .IN1(n7273), .IN2(n3636), .QN(N4376) );
  INVX0 U7982 ( .INP(n4479), .ZN(n7273) );
  NOR2X0 U7983 ( .IN1(n7274), .IN2(n3637), .QN(N4375) );
  INVX0 U7984 ( .INP(n4478), .ZN(n7274) );
  NOR2X0 U7985 ( .IN1(n7275), .IN2(n3638), .QN(N4374) );
  NOR2X0 U7986 ( .IN1(n7276), .IN2(n3639), .QN(N4373) );
  NOR2X0 U7987 ( .IN1(n7277), .IN2(n3640), .QN(N4372) );
  NOR2X0 U7988 ( .IN1(n7278), .IN2(n3641), .QN(N4371) );
  NOR2X0 U7989 ( .IN1(n7279), .IN2(n3642), .QN(N4370) );
  MUX21X1 U7990 ( .IN1(N325), .IN2(n9119), .S(n9191), .Q(N437) );
  NOR2X0 U7991 ( .IN1(n7280), .IN2(n3643), .QN(N4369) );
  NOR2X0 U7992 ( .IN1(n7281), .IN2(n3644), .QN(N4368) );
  NOR2X0 U7993 ( .IN1(n7282), .IN2(n3645), .QN(N4367) );
  NOR2X0 U7994 ( .IN1(n7283), .IN2(n3646), .QN(N4366) );
  NOR2X0 U7995 ( .IN1(n7284), .IN2(n3647), .QN(N4365) );
  NOR2X0 U7996 ( .IN1(n7285), .IN2(n3648), .QN(N4364) );
  NOR2X0 U7997 ( .IN1(n7286), .IN2(n3649), .QN(N4363) );
  NOR2X0 U7998 ( .IN1(n7287), .IN2(n3650), .QN(N4362) );
  NOR2X0 U7999 ( .IN1(n7288), .IN2(n3651), .QN(N4361) );
  NOR2X0 U8000 ( .IN1(n7289), .IN2(n3652), .QN(N4360) );
  MUX21X1 U8001 ( .IN1(N324), .IN2(n9121), .S(n9191), .Q(N436) );
  NOR2X0 U8002 ( .IN1(n7290), .IN2(n3653), .QN(N4359) );
  NOR2X0 U8003 ( .IN1(n7291), .IN2(n3654), .QN(N4358) );
  NOR2X0 U8004 ( .IN1(n7292), .IN2(n3655), .QN(N4357) );
  NOR2X0 U8005 ( .IN1(n7293), .IN2(n3656), .QN(N4356) );
  NOR2X0 U8006 ( .IN1(n7294), .IN2(n3657), .QN(N4355) );
  NOR2X0 U8007 ( .IN1(n7295), .IN2(n3658), .QN(N4354) );
  NOR2X0 U8008 ( .IN1(n7296), .IN2(n3659), .QN(N4353) );
  NOR2X0 U8009 ( .IN1(n7297), .IN2(n3660), .QN(N4352) );
  NOR2X0 U8010 ( .IN1(n7298), .IN2(n3661), .QN(N4351) );
  MUX21X1 U8011 ( .IN1(N323), .IN2(n9122), .S(n9191), .Q(N435) );
  AO221X1 U8012 ( .IN1(n8051), .IN2(n7232), .IN3(n7583), .IN4(n8052), .IN5(
        n7584), .Q(N4140) );
  OR2X1 U8013 ( .IN1(n8053), .IN2(n8054), .Q(n8051) );
  AO221X1 U8014 ( .IN1(n7581), .IN2(n8052), .IN3(n7583), .IN4(n8055), .IN5(
        n7584), .Q(N4139) );
  AO221X1 U8015 ( .IN1(n7581), .IN2(n8055), .IN3(n7583), .IN4(n8056), .IN5(
        n7584), .Q(N4138) );
  AO221X1 U8016 ( .IN1(n7581), .IN2(n8056), .IN3(n7583), .IN4(n8057), .IN5(
        n7584), .Q(N4137) );
  AO222X1 U8017 ( .IN1(n7623), .IN2(n8055), .IN3(n8052), .IN4(n7626), .IN5(
        n7625), .IN6(n8058), .Q(n8056) );
  AO221X1 U8018 ( .IN1(n7581), .IN2(n8057), .IN3(n7583), .IN4(n8059), .IN5(
        n7584), .Q(N4136) );
  AO222X1 U8019 ( .IN1(n7623), .IN2(n8058), .IN3(n8055), .IN4(n7626), .IN5(
        n7625), .IN6(n8060), .Q(n8057) );
  AO222X1 U8020 ( .IN1(n7631), .IN2(n8061), .IN3(n8052), .IN4(n7629), .IN5(
        n7633), .IN6(n7232), .Q(n8055) );
  AO221X1 U8021 ( .IN1(n7581), .IN2(n8059), .IN3(n7583), .IN4(n8062), .IN5(
        n7584), .Q(N4135) );
  AO222X1 U8022 ( .IN1(n7623), .IN2(n8060), .IN3(n8058), .IN4(n7626), .IN5(
        n7625), .IN6(n8063), .Q(n8059) );
  AO222X1 U8023 ( .IN1(n7629), .IN2(n8061), .IN3(n7633), .IN4(n8052), .IN5(
        n7631), .IN6(n8064), .Q(n8058) );
  AO221X1 U8024 ( .IN1(n7581), .IN2(n8062), .IN3(n7583), .IN4(n8065), .IN5(
        n7584), .Q(N4134) );
  AO222X1 U8025 ( .IN1(n7623), .IN2(n8063), .IN3(n8060), .IN4(n7626), .IN5(
        n7625), .IN6(n8066), .Q(n8062) );
  AO222X1 U8026 ( .IN1(n7629), .IN2(n8064), .IN3(n7633), .IN4(n8061), .IN5(
        n7631), .IN6(n8067), .Q(n8060) );
  AO222X1 U8027 ( .IN1(n7637), .IN2(n8068), .IN3(n8052), .IN4(n7635), .IN5(
        n7638), .IN6(n7232), .Q(n8061) );
  AO221X1 U8028 ( .IN1(n7581), .IN2(n8065), .IN3(n7583), .IN4(n8069), .IN5(
        n7584), .Q(N4133) );
  AO222X1 U8029 ( .IN1(n7623), .IN2(n8066), .IN3(n8063), .IN4(n7626), .IN5(
        n7625), .IN6(n8070), .Q(n8065) );
  AO222X1 U8030 ( .IN1(n7629), .IN2(n8067), .IN3(n7633), .IN4(n8064), .IN5(
        n7631), .IN6(n8071), .Q(n8063) );
  AO222X1 U8031 ( .IN1(n7635), .IN2(n8068), .IN3(n8052), .IN4(n7638), .IN5(
        n7637), .IN6(n8072), .Q(n8064) );
  MUX21X1 U8032 ( .IN1(n8073), .IN2(n7232), .S(n7666), .Q(n8052) );
  AO221X1 U8033 ( .IN1(n7581), .IN2(n8069), .IN3(n7583), .IN4(n8074), .IN5(
        n7584), .Q(N4132) );
  AO222X1 U8034 ( .IN1(n7623), .IN2(n8070), .IN3(n8066), .IN4(n7626), .IN5(
        n7625), .IN6(n8075), .Q(n8069) );
  AO222X1 U8035 ( .IN1(n7629), .IN2(n8071), .IN3(n7633), .IN4(n8067), .IN5(
        n7631), .IN6(n8076), .Q(n8066) );
  AO222X1 U8036 ( .IN1(n7635), .IN2(n8072), .IN3(n8068), .IN4(n7638), .IN5(
        n7637), .IN6(n8077), .Q(n8067) );
  AO222X1 U8037 ( .IN1(n8078), .IN2(n8079), .IN3(n8073), .IN4(n7659), .IN5(
        n7660), .IN6(n7232), .Q(n8068) );
  AO221X1 U8038 ( .IN1(n7581), .IN2(n8074), .IN3(n7583), .IN4(n8080), .IN5(
        n7584), .Q(N4131) );
  AO221X1 U8039 ( .IN1(n7581), .IN2(n8080), .IN3(n7583), .IN4(n8081), .IN5(
        n7584), .Q(N4130) );
  AO221X1 U8040 ( .IN1(n7581), .IN2(n8081), .IN3(n7583), .IN4(n8082), .IN5(
        n7584), .Q(N4129) );
  AO222X1 U8041 ( .IN1(n7598), .IN2(n8080), .IN3(n8074), .IN4(n7599), .IN5(
        n8083), .IN6(n8084), .Q(n8081) );
  AO222X1 U8042 ( .IN1(n7623), .IN2(n8075), .IN3(n8070), .IN4(n7626), .IN5(
        n7625), .IN6(n8085), .Q(n8074) );
  AO222X1 U8043 ( .IN1(n7629), .IN2(n8076), .IN3(n7633), .IN4(n8071), .IN5(
        n7631), .IN6(n8086), .Q(n8070) );
  AO222X1 U8044 ( .IN1(n7635), .IN2(n8077), .IN3(n8072), .IN4(n7638), .IN5(
        n7637), .IN6(n8087), .Q(n8071) );
  AO221X1 U8045 ( .IN1(n7581), .IN2(n8082), .IN3(n7583), .IN4(n8088), .IN5(
        n7584), .Q(N4128) );
  AO221X1 U8046 ( .IN1(n7581), .IN2(n8088), .IN3(n7583), .IN4(n8089), .IN5(
        n7584), .Q(N4127) );
  AO221X1 U8047 ( .IN1(n7581), .IN2(n8089), .IN3(n7583), .IN4(n8090), .IN5(
        n7584), .Q(N4126) );
  AO222X1 U8048 ( .IN1(n7592), .IN2(n8088), .IN3(n7596), .IN4(n8082), .IN5(
        n7594), .IN6(n8091), .Q(n8089) );
  AO222X1 U8049 ( .IN1(n7598), .IN2(n8084), .IN3(n8080), .IN4(n7599), .IN5(
        n8083), .IN6(n8092), .Q(n8082) );
  AO221X1 U8050 ( .IN1(n7581), .IN2(n8090), .IN3(n7583), .IN4(n8093), .IN5(
        n7584), .Q(N4125) );
  AO222X1 U8051 ( .IN1(n7592), .IN2(n8091), .IN3(n7596), .IN4(n8088), .IN5(
        n7594), .IN6(n8094), .Q(n8090) );
  AO222X1 U8052 ( .IN1(n7598), .IN2(n8092), .IN3(n8084), .IN4(n7599), .IN5(
        n8083), .IN6(n8095), .Q(n8088) );
  AO221X1 U8053 ( .IN1(n7581), .IN2(n8093), .IN3(n7583), .IN4(n8096), .IN5(
        n7584), .Q(N4124) );
  AO222X1 U8054 ( .IN1(n7592), .IN2(n8094), .IN3(n7596), .IN4(n8091), .IN5(
        n7594), .IN6(n8097), .Q(n8093) );
  AO222X1 U8055 ( .IN1(n7598), .IN2(n8095), .IN3(n8092), .IN4(n7599), .IN5(
        n8083), .IN6(n8098), .Q(n8091) );
  AO222X1 U8056 ( .IN1(n7609), .IN2(n8084), .IN3(n8080), .IN4(n7606), .IN5(
        n8099), .IN6(n8100), .Q(n8092) );
  AO222X1 U8057 ( .IN1(n7623), .IN2(n8085), .IN3(n8075), .IN4(n7626), .IN5(
        n7625), .IN6(n8101), .Q(n8080) );
  AO222X1 U8058 ( .IN1(n7629), .IN2(n8086), .IN3(n7633), .IN4(n8076), .IN5(
        n7631), .IN6(n8102), .Q(n8075) );
  AO222X1 U8059 ( .IN1(n7635), .IN2(n8087), .IN3(n8077), .IN4(n7638), .IN5(
        n7637), .IN6(n8103), .Q(n8076) );
  AO221X1 U8060 ( .IN1(n7581), .IN2(n8096), .IN3(n7583), .IN4(n8104), .IN5(
        n7584), .Q(N4123) );
  AO222X1 U8061 ( .IN1(n7592), .IN2(n8097), .IN3(n7596), .IN4(n8094), .IN5(
        n7594), .IN6(n8105), .Q(n8096) );
  AO222X1 U8062 ( .IN1(n7598), .IN2(n8098), .IN3(n8095), .IN4(n7599), .IN5(
        n8083), .IN6(n8106), .Q(n8094) );
  AO222X1 U8063 ( .IN1(n7609), .IN2(n8100), .IN3(n8084), .IN4(n7606), .IN5(
        n8099), .IN6(n8107), .Q(n8095) );
  AO221X1 U8064 ( .IN1(n7581), .IN2(n8104), .IN3(n7583), .IN4(n8108), .IN5(
        n7584), .Q(N4122) );
  AO221X1 U8065 ( .IN1(n7581), .IN2(n8108), .IN3(n7583), .IN4(n8109), .IN5(
        n7584), .Q(N4121) );
  AO221X1 U8066 ( .IN1(n7581), .IN2(n8109), .IN3(n7583), .IN4(n8110), .IN5(
        n7584), .Q(N4120) );
  AO222X1 U8067 ( .IN1(n7586), .IN2(n8108), .IN3(n7590), .IN4(n8104), .IN5(
        n7588), .IN6(n8111), .Q(n8109) );
  AO222X1 U8068 ( .IN1(n7592), .IN2(n8105), .IN3(n7596), .IN4(n8097), .IN5(
        n7594), .IN6(n8112), .Q(n8104) );
  AO222X1 U8069 ( .IN1(n7598), .IN2(n8106), .IN3(n8098), .IN4(n7599), .IN5(
        n8083), .IN6(n8113), .Q(n8097) );
  AO222X1 U8070 ( .IN1(n7609), .IN2(n8107), .IN3(n8100), .IN4(n7606), .IN5(
        n8099), .IN6(n8114), .Q(n8098) );
  AO221X1 U8071 ( .IN1(n7581), .IN2(n8110), .IN3(n7583), .IN4(n8115), .IN5(
        n7584), .Q(N4119) );
  AO222X1 U8072 ( .IN1(n7586), .IN2(n8111), .IN3(n7590), .IN4(n8108), .IN5(
        n7588), .IN6(n8116), .Q(n8110) );
  AO222X1 U8073 ( .IN1(n7592), .IN2(n8112), .IN3(n7596), .IN4(n8105), .IN5(
        n7594), .IN6(n8117), .Q(n8108) );
  AO222X1 U8074 ( .IN1(n7598), .IN2(n8113), .IN3(n8106), .IN4(n7599), .IN5(
        n8083), .IN6(n8118), .Q(n8105) );
  AO222X1 U8075 ( .IN1(n7609), .IN2(n8114), .IN3(n8107), .IN4(n7606), .IN5(
        n8099), .IN6(n8119), .Q(n8106) );
  AO222X1 U8076 ( .IN1(n7611), .IN2(n8100), .IN3(n7615), .IN4(n8084), .IN5(
        n7613), .IN6(n8120), .Q(n8107) );
  AO222X1 U8077 ( .IN1(n7623), .IN2(n8101), .IN3(n8085), .IN4(n7626), .IN5(
        n7625), .IN6(n8121), .Q(n8084) );
  AO222X1 U8078 ( .IN1(n7629), .IN2(n8102), .IN3(n7633), .IN4(n8086), .IN5(
        n7631), .IN6(n8122), .Q(n8085) );
  AO222X1 U8079 ( .IN1(n7635), .IN2(n8103), .IN3(n8087), .IN4(n7638), .IN5(
        n7637), .IN6(n8123), .Q(n8086) );
  AO222X1 U8080 ( .IN1(n7641), .IN2(n8087), .IN3(n8077), .IN4(n7644), .IN5(
        n7643), .IN6(n8124), .Q(n8103) );
  AO221X1 U8081 ( .IN1(n7581), .IN2(n8115), .IN3(n7583), .IN4(n8125), .IN5(
        n7584), .Q(N4118) );
  AO222X1 U8082 ( .IN1(n7586), .IN2(n8116), .IN3(n7590), .IN4(n8111), .IN5(
        n7588), .IN6(n8126), .Q(n8115) );
  AO222X1 U8083 ( .IN1(n7592), .IN2(n8117), .IN3(n7596), .IN4(n8112), .IN5(
        n7594), .IN6(n8127), .Q(n8111) );
  AO222X1 U8084 ( .IN1(n7598), .IN2(n8118), .IN3(n8113), .IN4(n7599), .IN5(
        n8083), .IN6(n8128), .Q(n8112) );
  AO222X1 U8085 ( .IN1(n7609), .IN2(n8119), .IN3(n8114), .IN4(n7606), .IN5(
        n8099), .IN6(n8129), .Q(n8113) );
  AO222X1 U8086 ( .IN1(n7611), .IN2(n8120), .IN3(n7615), .IN4(n8100), .IN5(
        n7613), .IN6(n8130), .Q(n8114) );
  AO222X1 U8087 ( .IN1(n7623), .IN2(n8121), .IN3(n8101), .IN4(n7626), .IN5(
        n7625), .IN6(n8131), .Q(n8100) );
  AO222X1 U8088 ( .IN1(n7629), .IN2(n8122), .IN3(n7633), .IN4(n8102), .IN5(
        n7631), .IN6(n8132), .Q(n8101) );
  AO221X1 U8089 ( .IN1(n7581), .IN2(n8125), .IN3(n7583), .IN4(n8133), .IN5(
        n7584), .Q(N4117) );
  AO222X1 U8090 ( .IN1(n7586), .IN2(n8126), .IN3(n7590), .IN4(n8116), .IN5(
        n7588), .IN6(n8134), .Q(n8125) );
  AO222X1 U8091 ( .IN1(n7592), .IN2(n8127), .IN3(n7596), .IN4(n8117), .IN5(
        n7594), .IN6(n8135), .Q(n8116) );
  AO222X1 U8092 ( .IN1(n7598), .IN2(n8128), .IN3(n8118), .IN4(n7599), .IN5(
        n8083), .IN6(n8136), .Q(n8117) );
  AO222X1 U8093 ( .IN1(n7609), .IN2(n8129), .IN3(n8119), .IN4(n7606), .IN5(
        n8099), .IN6(n8137), .Q(n8118) );
  AO222X1 U8094 ( .IN1(n7611), .IN2(n8130), .IN3(n7615), .IN4(n8120), .IN5(
        n7613), .IN6(n8138), .Q(n8119) );
  AO222X1 U8095 ( .IN1(n7623), .IN2(n8131), .IN3(n8121), .IN4(n7626), .IN5(
        n7625), .IN6(n8139), .Q(n8120) );
  AO222X1 U8096 ( .IN1(n7629), .IN2(n8132), .IN3(n7633), .IN4(n8122), .IN5(
        n7631), .IN6(n8140), .Q(n8121) );
  AO222X1 U8097 ( .IN1(n7635), .IN2(n8102), .IN3(n8123), .IN4(n7638), .IN5(
        n7637), .IN6(n8141), .Q(n8122) );
  AO222X1 U8098 ( .IN1(n7641), .IN2(n8124), .IN3(n8087), .IN4(n7644), .IN5(
        n7643), .IN6(n8142), .Q(n8123) );
  AO222X1 U8099 ( .IN1(n7647), .IN2(n8077), .IN3(n8072), .IN4(n7650), .IN5(
        n7649), .IN6(n8143), .Q(n8087) );
  AO222X1 U8100 ( .IN1(n7659), .IN2(n8079), .IN3(n8073), .IN4(n7660), .IN5(
        n8078), .IN6(n8144), .Q(n8072) );
  MUX21X1 U8101 ( .IN1(n7232), .IN2(n8145), .S(n8146), .Q(n8073) );
  AO221X1 U8102 ( .IN1(n7581), .IN2(n8133), .IN3(n7583), .IN4(n8147), .IN5(
        n7584), .Q(N4116) );
  AO222X1 U8103 ( .IN1(n7586), .IN2(n8134), .IN3(n7590), .IN4(n8126), .IN5(
        n7588), .IN6(n8148), .Q(n8133) );
  AO222X1 U8104 ( .IN1(n7592), .IN2(n8135), .IN3(n7596), .IN4(n8127), .IN5(
        n7594), .IN6(n8149), .Q(n8126) );
  AO222X1 U8105 ( .IN1(n7598), .IN2(n8136), .IN3(n8128), .IN4(n7599), .IN5(
        n8083), .IN6(n8150), .Q(n8127) );
  AO222X1 U8106 ( .IN1(n7609), .IN2(n8137), .IN3(n8129), .IN4(n7606), .IN5(
        n8099), .IN6(n8151), .Q(n8128) );
  AO222X1 U8107 ( .IN1(n7611), .IN2(n8138), .IN3(n7615), .IN4(n8130), .IN5(
        n7613), .IN6(n8152), .Q(n8129) );
  AO222X1 U8108 ( .IN1(n7623), .IN2(n8139), .IN3(n8131), .IN4(n7626), .IN5(
        n7625), .IN6(n8153), .Q(n8130) );
  AO222X1 U8109 ( .IN1(n7629), .IN2(n8140), .IN3(n7633), .IN4(n8132), .IN5(
        n7631), .IN6(n8154), .Q(n8131) );
  AO222X1 U8110 ( .IN1(n7635), .IN2(n8141), .IN3(n8102), .IN4(n7638), .IN5(
        n7637), .IN6(n8155), .Q(n8132) );
  AO222X1 U8111 ( .IN1(n7641), .IN2(n8142), .IN3(n8124), .IN4(n7644), .IN5(
        n7643), .IN6(n8156), .Q(n8102) );
  AO222X1 U8112 ( .IN1(n7647), .IN2(n8143), .IN3(n8077), .IN4(n7650), .IN5(
        n7649), .IN6(n8157), .Q(n8124) );
  AO222X1 U8113 ( .IN1(n8078), .IN2(n8158), .IN3(n8079), .IN4(n7660), .IN5(
        n7659), .IN6(n8144), .Q(n8077) );
  AO222X1 U8114 ( .IN1(n8145), .IN2(n7670), .IN3(n8146), .IN4(n8159), .IN5(
        n7668), .IN6(n7232), .Q(n8079) );
  AO221X1 U8115 ( .IN1(n7581), .IN2(n8147), .IN3(n7583), .IN4(n8160), .IN5(
        n7584), .Q(N4115) );
  AO222X1 U8116 ( .IN1(n7586), .IN2(n8148), .IN3(n7590), .IN4(n8134), .IN5(
        n7588), .IN6(n8161), .Q(n8147) );
  AO222X1 U8117 ( .IN1(n7592), .IN2(n8149), .IN3(n7596), .IN4(n8135), .IN5(
        n7594), .IN6(n8162), .Q(n8134) );
  AO222X1 U8118 ( .IN1(n7598), .IN2(n8150), .IN3(n8136), .IN4(n7599), .IN5(
        n8083), .IN6(n8163), .Q(n8135) );
  AO222X1 U8119 ( .IN1(n7609), .IN2(n8151), .IN3(n8137), .IN4(n7606), .IN5(
        n8099), .IN6(n8164), .Q(n8136) );
  AO222X1 U8120 ( .IN1(n7611), .IN2(n8152), .IN3(n7615), .IN4(n8138), .IN5(
        n7613), .IN6(n8165), .Q(n8137) );
  AO221X1 U8121 ( .IN1(n7581), .IN2(n8160), .IN3(n7583), .IN4(n8166), .IN5(
        n7584), .Q(N4114) );
  AO222X1 U8122 ( .IN1(n7586), .IN2(n8161), .IN3(n7590), .IN4(n8148), .IN5(
        n7588), .IN6(n8167), .Q(n8160) );
  AO222X1 U8123 ( .IN1(n7592), .IN2(n8162), .IN3(n7596), .IN4(n8149), .IN5(
        n7594), .IN6(n8168), .Q(n8148) );
  AO222X1 U8124 ( .IN1(n7598), .IN2(n8163), .IN3(n8150), .IN4(n7599), .IN5(
        n8083), .IN6(n8169), .Q(n8149) );
  AO222X1 U8125 ( .IN1(n7609), .IN2(n8164), .IN3(n8151), .IN4(n7606), .IN5(
        n8099), .IN6(n8170), .Q(n8150) );
  AO222X1 U8126 ( .IN1(n7611), .IN2(n8165), .IN3(n7615), .IN4(n8152), .IN5(
        n7613), .IN6(n8171), .Q(n8151) );
  AO221X1 U8127 ( .IN1(n7581), .IN2(n8166), .IN3(n7583), .IN4(n8172), .IN5(
        n7584), .Q(N4113) );
  AO222X1 U8128 ( .IN1(n7586), .IN2(n8167), .IN3(n7590), .IN4(n8161), .IN5(
        n7588), .IN6(n8173), .Q(n8166) );
  AO222X1 U8129 ( .IN1(n7592), .IN2(n8168), .IN3(n7596), .IN4(n8162), .IN5(
        n7594), .IN6(n8174), .Q(n8161) );
  AO222X1 U8130 ( .IN1(n7598), .IN2(n8169), .IN3(n8163), .IN4(n7599), .IN5(
        n8083), .IN6(n8175), .Q(n8162) );
  AO222X1 U8131 ( .IN1(n7609), .IN2(n8170), .IN3(n8164), .IN4(n7606), .IN5(
        n8099), .IN6(n8176), .Q(n8163) );
  AO222X1 U8132 ( .IN1(n7611), .IN2(n8171), .IN3(n7615), .IN4(n8165), .IN5(
        n7613), .IN6(n8177), .Q(n8164) );
  AO222X1 U8133 ( .IN1(n7617), .IN2(n8152), .IN3(n7621), .IN4(n8138), .IN5(
        n7619), .IN6(n8178), .Q(n8165) );
  AO222X1 U8134 ( .IN1(n7623), .IN2(n8153), .IN3(n8139), .IN4(n7626), .IN5(
        n7625), .IN6(n8179), .Q(n8138) );
  AO222X1 U8135 ( .IN1(n7629), .IN2(n8154), .IN3(n7633), .IN4(n8140), .IN5(
        n7631), .IN6(n8180), .Q(n8139) );
  AO222X1 U8136 ( .IN1(n7635), .IN2(n8155), .IN3(n8141), .IN4(n7638), .IN5(
        n7637), .IN6(n8181), .Q(n8140) );
  AO222X1 U8137 ( .IN1(n7641), .IN2(n8156), .IN3(n8142), .IN4(n7644), .IN5(
        n7643), .IN6(n8182), .Q(n8141) );
  AO222X1 U8138 ( .IN1(n7647), .IN2(n8157), .IN3(n8143), .IN4(n7650), .IN5(
        n7649), .IN6(n8183), .Q(n8142) );
  AO221X1 U8139 ( .IN1(n7581), .IN2(n8172), .IN3(n7583), .IN4(n8184), .IN5(
        n7584), .Q(N4112) );
  AO222X1 U8140 ( .IN1(n7588), .IN2(n8185), .IN3(n7590), .IN4(n8167), .IN5(
        n7586), .IN6(n8173), .Q(n8172) );
  AO222X1 U8141 ( .IN1(n7594), .IN2(n8186), .IN3(n7596), .IN4(n8168), .IN5(
        n7592), .IN6(n8174), .Q(n8167) );
  AO222X1 U8142 ( .IN1(n8083), .IN2(n8187), .IN3(n8169), .IN4(n7599), .IN5(
        n7598), .IN6(n8175), .Q(n8168) );
  AO222X1 U8143 ( .IN1(n8099), .IN2(n8188), .IN3(n8170), .IN4(n7606), .IN5(
        n7609), .IN6(n8176), .Q(n8169) );
  AO222X1 U8144 ( .IN1(n7613), .IN2(n8189), .IN3(n7615), .IN4(n8171), .IN5(
        n7611), .IN6(n8177), .Q(n8170) );
  AO222X1 U8145 ( .IN1(n7619), .IN2(n8190), .IN3(n7621), .IN4(n8152), .IN5(
        n7617), .IN6(n8178), .Q(n8171) );
  AO222X1 U8146 ( .IN1(n7625), .IN2(n8191), .IN3(n8153), .IN4(n7626), .IN5(
        n7623), .IN6(n8179), .Q(n8152) );
  AO222X1 U8147 ( .IN1(n7631), .IN2(n8192), .IN3(n7633), .IN4(n8154), .IN5(
        n7629), .IN6(n8180), .Q(n8153) );
  AO222X1 U8148 ( .IN1(n7637), .IN2(n8193), .IN3(n8155), .IN4(n7638), .IN5(
        n7635), .IN6(n8181), .Q(n8154) );
  AO222X1 U8149 ( .IN1(n7643), .IN2(n8194), .IN3(n8156), .IN4(n7644), .IN5(
        n7641), .IN6(n8182), .Q(n8155) );
  AO222X1 U8150 ( .IN1(n7649), .IN2(n8195), .IN3(n8157), .IN4(n7650), .IN5(
        n7647), .IN6(n8183), .Q(n8156) );
  AO221X1 U8151 ( .IN1(n7583), .IN2(n8196), .IN3(n7581), .IN4(n8184), .IN5(
        n7584), .Q(N4111) );
  AO222X1 U8152 ( .IN1(n7590), .IN2(n8173), .IN3(n7586), .IN4(n8185), .IN5(
        n7588), .IN6(n8197), .Q(n8184) );
  AO222X1 U8153 ( .IN1(n7596), .IN2(n8174), .IN3(n7592), .IN4(n8186), .IN5(
        n7594), .IN6(n8198), .Q(n8173) );
  AO222X1 U8154 ( .IN1(n8175), .IN2(n7599), .IN3(n7598), .IN4(n8187), .IN5(
        n8083), .IN6(n8199), .Q(n8174) );
  AO222X1 U8155 ( .IN1(n8176), .IN2(n7606), .IN3(n7609), .IN4(n8188), .IN5(
        n8099), .IN6(n8200), .Q(n8175) );
  AO222X1 U8156 ( .IN1(n7615), .IN2(n8177), .IN3(n7611), .IN4(n8189), .IN5(
        n7613), .IN6(n8201), .Q(n8176) );
  AO222X1 U8157 ( .IN1(n7621), .IN2(n8178), .IN3(n7617), .IN4(n8190), .IN5(
        n7619), .IN6(n8202), .Q(n8177) );
  AO222X1 U8158 ( .IN1(n8179), .IN2(n7626), .IN3(n7623), .IN4(n8191), .IN5(
        n7625), .IN6(n8203), .Q(n8178) );
  AO222X1 U8159 ( .IN1(n7633), .IN2(n8180), .IN3(n7629), .IN4(n8192), .IN5(
        n7631), .IN6(n8204), .Q(n8179) );
  AO222X1 U8160 ( .IN1(n8181), .IN2(n7638), .IN3(n7635), .IN4(n8193), .IN5(
        n7637), .IN6(n8205), .Q(n8180) );
  AO222X1 U8161 ( .IN1(n8182), .IN2(n7644), .IN3(n7641), .IN4(n8194), .IN5(
        n7643), .IN6(n8206), .Q(n8181) );
  AO222X1 U8162 ( .IN1(n8183), .IN2(n7650), .IN3(n7647), .IN4(n8195), .IN5(
        n7649), .IN6(n8207), .Q(n8182) );
  AO222X1 U8163 ( .IN1(n7657), .IN2(n8143), .IN3(n7653), .IN4(n8157), .IN5(
        n7655), .IN6(n8208), .Q(n8183) );
  AO222X1 U8164 ( .IN1(n8144), .IN2(n7660), .IN3(n7659), .IN4(n8158), .IN5(
        n8078), .IN6(n8209), .Q(n8143) );
  AO222X1 U8165 ( .IN1(n7668), .IN2(n8145), .IN3(n7670), .IN4(n8159), .IN5(
        n8146), .IN6(n8210), .Q(n8144) );
  MUX21X1 U8166 ( .IN1(n7233), .IN2(n7232), .S(n8211), .Q(n8145) );
  AO221X1 U8167 ( .IN1(n7581), .IN2(n8196), .IN3(n7583), .IN4(n7580), .IN5(
        n7584), .Q(N4110) );
  NOR2X0 U8168 ( .IN1(n7528), .IN2(n3661), .QN(n7584) );
  AO222X1 U8169 ( .IN1(n7588), .IN2(n7585), .IN3(n7586), .IN4(n7589), .IN5(
        n7590), .IN6(n8197), .Q(n7580) );
  AO222X1 U8170 ( .IN1(n7594), .IN2(n7591), .IN3(n7592), .IN4(n7595), .IN5(
        n7596), .IN6(n8212), .Q(n7585) );
  AO222X1 U8171 ( .IN1(n8083), .IN2(n7597), .IN3(n7598), .IN4(n7600), .IN5(
        n8213), .IN6(n7599), .Q(n7591) );
  AO222X1 U8172 ( .IN1(n8099), .IN2(n7608), .IN3(n7609), .IN4(n7607), .IN5(
        n8214), .IN6(n7606), .Q(n7597) );
  AO222X1 U8173 ( .IN1(n7613), .IN2(n7610), .IN3(n7611), .IN4(n7614), .IN5(
        n7615), .IN6(n8215), .Q(n7608) );
  AO222X1 U8174 ( .IN1(n7619), .IN2(n7616), .IN3(n7617), .IN4(n7620), .IN5(
        n7621), .IN6(n8216), .Q(n7610) );
  AO222X1 U8175 ( .IN1(n7625), .IN2(n7622), .IN3(n7623), .IN4(n7627), .IN5(
        n8217), .IN6(n7626), .Q(n7616) );
  AO222X1 U8176 ( .IN1(n7631), .IN2(n7628), .IN3(n7629), .IN4(n7632), .IN5(
        n7633), .IN6(n8218), .Q(n7622) );
  AO222X1 U8177 ( .IN1(n7637), .IN2(n7634), .IN3(n7635), .IN4(n7639), .IN5(
        n8219), .IN6(n7638), .Q(n7628) );
  AO222X1 U8178 ( .IN1(n7643), .IN2(n7640), .IN3(n7641), .IN4(n7645), .IN5(
        n8220), .IN6(n7644), .Q(n7634) );
  AO222X1 U8179 ( .IN1(n7649), .IN2(n7646), .IN3(n7647), .IN4(n7651), .IN5(
        n8221), .IN6(n7650), .Q(n7640) );
  AO222X1 U8180 ( .IN1(n7655), .IN2(n7652), .IN3(n7653), .IN4(n7656), .IN5(
        n7657), .IN6(n8222), .Q(n7646) );
  AO222X1 U8181 ( .IN1(n8078), .IN2(n7658), .IN3(n7659), .IN4(n7661), .IN5(
        n8223), .IN6(n7660), .Q(n7652) );
  AO222X1 U8182 ( .IN1(n8146), .IN2(n7669), .IN3(n7670), .IN4(n7667), .IN5(
        n7668), .IN6(n8224), .Q(n7658) );
  AO222X1 U8183 ( .IN1(n7672), .IN2(n7262), .IN3(n7671), .IN4(n7261), .IN5(
        n8225), .IN6(n7263), .Q(n7669) );
  INVX0 U8184 ( .INP(n3630), .ZN(n7263) );
  NOR3X0 U8185 ( .IN1(n8053), .IN2(n8054), .IN3(n8049), .QN(n7583) );
  AO222X1 U8186 ( .IN1(n7590), .IN2(n8185), .IN3(n7588), .IN4(n7589), .IN5(
        n7586), .IN6(n8197), .Q(n8196) );
  AO222X1 U8187 ( .IN1(n7596), .IN2(n8198), .IN3(n7592), .IN4(n8226), .IN5(
        n7594), .IN6(n8212), .Q(n8197) );
  XOR2X1 U8188 ( .IN1(n7712), .IN2(n8227), .Q(n7586) );
  AO222X1 U8189 ( .IN1(n7596), .IN2(n8226), .IN3(n7594), .IN4(n7595), .IN5(
        n7592), .IN6(n8212), .Q(n7589) );
  AO222X1 U8190 ( .IN1(n8228), .IN2(n7599), .IN3(n7598), .IN4(n8229), .IN5(
        n8083), .IN6(n8213), .Q(n8212) );
  AO222X1 U8191 ( .IN1(n8229), .IN2(n7599), .IN3(n8083), .IN4(n7600), .IN5(
        n7598), .IN6(n8213), .Q(n7595) );
  AO222X1 U8192 ( .IN1(n8230), .IN2(n7606), .IN3(n7609), .IN4(n8231), .IN5(
        n8099), .IN6(n8214), .Q(n8213) );
  AO222X1 U8193 ( .IN1(n8231), .IN2(n7606), .IN3(n8099), .IN4(n7607), .IN5(
        n7609), .IN6(n8214), .Q(n7600) );
  AO222X1 U8194 ( .IN1(n7615), .IN2(n8232), .IN3(n7611), .IN4(n8233), .IN5(
        n7613), .IN6(n8215), .Q(n8214) );
  AO222X1 U8195 ( .IN1(n7615), .IN2(n8233), .IN3(n7613), .IN4(n7614), .IN5(
        n7611), .IN6(n8215), .Q(n7607) );
  AO222X1 U8196 ( .IN1(n7621), .IN2(n8234), .IN3(n7617), .IN4(n8235), .IN5(
        n7619), .IN6(n8216), .Q(n8215) );
  AO222X1 U8197 ( .IN1(n7621), .IN2(n8235), .IN3(n7619), .IN4(n7620), .IN5(
        n7617), .IN6(n8216), .Q(n7614) );
  AO222X1 U8198 ( .IN1(n8236), .IN2(n7626), .IN3(n7623), .IN4(n8237), .IN5(
        n7625), .IN6(n8217), .Q(n8216) );
  AO222X1 U8199 ( .IN1(n8237), .IN2(n7626), .IN3(n7625), .IN4(n7627), .IN5(
        n7623), .IN6(n8217), .Q(n7620) );
  AO222X1 U8200 ( .IN1(n7631), .IN2(n8218), .IN3(n7629), .IN4(n8238), .IN5(
        n7633), .IN6(n8239), .Q(n8217) );
  AO222X1 U8201 ( .IN1(n7633), .IN2(n8238), .IN3(n7631), .IN4(n7632), .IN5(
        n7629), .IN6(n8218), .Q(n7627) );
  AO222X1 U8202 ( .IN1(n7637), .IN2(n8219), .IN3(n7635), .IN4(n8240), .IN5(
        n8241), .IN6(n7638), .Q(n8218) );
  AO222X1 U8203 ( .IN1(n8240), .IN2(n7638), .IN3(n7637), .IN4(n7639), .IN5(
        n7635), .IN6(n8219), .Q(n7632) );
  AO222X1 U8204 ( .IN1(n7643), .IN2(n8220), .IN3(n7641), .IN4(n8242), .IN5(
        n8243), .IN6(n7644), .Q(n8219) );
  AO222X1 U8205 ( .IN1(n8242), .IN2(n7644), .IN3(n7643), .IN4(n7645), .IN5(
        n7641), .IN6(n8220), .Q(n7639) );
  AO222X1 U8206 ( .IN1(n7649), .IN2(n8221), .IN3(n7647), .IN4(n8244), .IN5(
        n8245), .IN6(n7650), .Q(n8220) );
  AO222X1 U8207 ( .IN1(n8244), .IN2(n7650), .IN3(n7649), .IN4(n7651), .IN5(
        n7647), .IN6(n8221), .Q(n7645) );
  AO222X1 U8208 ( .IN1(n7655), .IN2(n8222), .IN3(n7653), .IN4(n8246), .IN5(
        n7657), .IN6(n8247), .Q(n8221) );
  AO222X1 U8209 ( .IN1(n7657), .IN2(n8246), .IN3(n7655), .IN4(n7656), .IN5(
        n7653), .IN6(n8222), .Q(n7651) );
  AO222X1 U8210 ( .IN1(n8078), .IN2(n8223), .IN3(n7659), .IN4(n8248), .IN5(
        n8249), .IN6(n7660), .Q(n8222) );
  AO222X1 U8211 ( .IN1(n8248), .IN2(n7660), .IN3(n8078), .IN4(n7661), .IN5(
        n7659), .IN6(n8223), .Q(n7656) );
  AO222X1 U8212 ( .IN1(n8146), .IN2(n8224), .IN3(n7670), .IN4(n8250), .IN5(
        n7668), .IN6(n8251), .Q(n8223) );
  AO222X1 U8213 ( .IN1(n7668), .IN2(n8250), .IN3(n8146), .IN4(n7667), .IN5(
        n7670), .IN6(n8224), .Q(n7661) );
  AO222X1 U8214 ( .IN1(n7672), .IN2(n7260), .IN3(n7671), .IN4(n7259), .IN5(
        n8225), .IN6(n7261), .Q(n8224) );
  AO222X1 U8215 ( .IN1(n7672), .IN2(n7261), .IN3(n7671), .IN4(n7260), .IN5(
        n8225), .IN6(n7262), .Q(n7667) );
  INVX0 U8216 ( .INP(n3631), .ZN(n7262) );
  INVX0 U8217 ( .INP(n3632), .ZN(n7261) );
  NOR2X0 U8218 ( .IN1(n7712), .IN2(n8227), .QN(n7588) );
  AO222X1 U8219 ( .IN1(n7594), .IN2(n8226), .IN3(n7596), .IN4(n8186), .IN5(
        n7592), .IN6(n8198), .Q(n8185) );
  AO222X1 U8220 ( .IN1(n8199), .IN2(n7599), .IN3(n7598), .IN4(n8252), .IN5(
        n8083), .IN6(n8228), .Q(n8198) );
  XOR2X1 U8221 ( .IN1(n8253), .IN2(n8254), .Q(n7592) );
  AO222X1 U8222 ( .IN1(n8083), .IN2(n8252), .IN3(n8187), .IN4(n7599), .IN5(
        n7598), .IN6(n8199), .Q(n8186) );
  AO222X1 U8223 ( .IN1(n8200), .IN2(n7606), .IN3(n7609), .IN4(n8255), .IN5(
        n8099), .IN6(n8256), .Q(n8199) );
  AO222X1 U8224 ( .IN1(n8099), .IN2(n8255), .IN3(n8188), .IN4(n7606), .IN5(
        n7609), .IN6(n8200), .Q(n8187) );
  AO222X1 U8225 ( .IN1(n7615), .IN2(n8201), .IN3(n7611), .IN4(n8257), .IN5(
        n7613), .IN6(n8258), .Q(n8200) );
  AO222X1 U8226 ( .IN1(n7613), .IN2(n8257), .IN3(n7615), .IN4(n8189), .IN5(
        n7611), .IN6(n8201), .Q(n8188) );
  AO222X1 U8227 ( .IN1(n7621), .IN2(n8202), .IN3(n7617), .IN4(n8259), .IN5(
        n7619), .IN6(n8260), .Q(n8201) );
  AO222X1 U8228 ( .IN1(n7619), .IN2(n8259), .IN3(n7621), .IN4(n8190), .IN5(
        n7617), .IN6(n8202), .Q(n8189) );
  AO222X1 U8229 ( .IN1(n8203), .IN2(n7626), .IN3(n7623), .IN4(n8261), .IN5(
        n7625), .IN6(n8262), .Q(n8202) );
  AO222X1 U8230 ( .IN1(n7625), .IN2(n8261), .IN3(n8191), .IN4(n7626), .IN5(
        n7623), .IN6(n8203), .Q(n8190) );
  AO222X1 U8231 ( .IN1(n7633), .IN2(n8204), .IN3(n7629), .IN4(n8263), .IN5(
        n7631), .IN6(n8264), .Q(n8203) );
  AO222X1 U8232 ( .IN1(n7631), .IN2(n8263), .IN3(n7633), .IN4(n8192), .IN5(
        n7629), .IN6(n8204), .Q(n8191) );
  AO222X1 U8233 ( .IN1(n8205), .IN2(n7638), .IN3(n7635), .IN4(n8265), .IN5(
        n7637), .IN6(n8266), .Q(n8204) );
  AO222X1 U8234 ( .IN1(n7637), .IN2(n8265), .IN3(n8193), .IN4(n7638), .IN5(
        n7635), .IN6(n8205), .Q(n8192) );
  AO222X1 U8235 ( .IN1(n8206), .IN2(n7644), .IN3(n7641), .IN4(n8267), .IN5(
        n7643), .IN6(n8268), .Q(n8205) );
  AO222X1 U8236 ( .IN1(n7643), .IN2(n8267), .IN3(n8194), .IN4(n7644), .IN5(
        n7641), .IN6(n8206), .Q(n8193) );
  AO222X1 U8237 ( .IN1(n8207), .IN2(n7650), .IN3(n7647), .IN4(n8269), .IN5(
        n7649), .IN6(n8270), .Q(n8206) );
  AO222X1 U8238 ( .IN1(n7649), .IN2(n8269), .IN3(n8195), .IN4(n7650), .IN5(
        n7647), .IN6(n8207), .Q(n8194) );
  AO222X1 U8239 ( .IN1(n7657), .IN2(n8208), .IN3(n7653), .IN4(n8271), .IN5(
        n7655), .IN6(n8272), .Q(n8207) );
  AO222X1 U8240 ( .IN1(n7655), .IN2(n8271), .IN3(n7657), .IN4(n8157), .IN5(
        n7653), .IN6(n8208), .Q(n8195) );
  AO222X1 U8241 ( .IN1(n8209), .IN2(n7660), .IN3(n7659), .IN4(n8273), .IN5(
        n8078), .IN6(n8274), .Q(n8208) );
  AO222X1 U8242 ( .IN1(n8078), .IN2(n8273), .IN3(n8158), .IN4(n7660), .IN5(
        n7659), .IN6(n8209), .Q(n8157) );
  AO222X1 U8243 ( .IN1(n7668), .IN2(n8210), .IN3(n7670), .IN4(n8275), .IN5(
        n8146), .IN6(n8276), .Q(n8209) );
  AO222X1 U8244 ( .IN1(n8146), .IN2(n8275), .IN3(n7668), .IN4(n8159), .IN5(
        n7670), .IN6(n8210), .Q(n8158) );
  AO222X1 U8245 ( .IN1(n7672), .IN2(n7234), .IN3(n7671), .IN4(n7233), .IN5(
        n8225), .IN6(n7235), .Q(n8210) );
  AO222X1 U8246 ( .IN1(n7672), .IN2(n7233), .IN3(n7671), .IN4(n7232), .IN5(
        n8225), .IN6(n7234), .Q(n8159) );
  INVX0 U8247 ( .INP(n3661), .ZN(n7232) );
  INVX0 U8248 ( .INP(n3660), .ZN(n7233) );
  AND2X1 U8249 ( .IN1(n8254), .IN2(n8253), .Q(n7596) );
  AO222X1 U8250 ( .IN1(n8083), .IN2(n8229), .IN3(n8252), .IN4(n7599), .IN5(
        n7598), .IN6(n8228), .Q(n8226) );
  AO222X1 U8251 ( .IN1(n8256), .IN2(n7606), .IN3(n7609), .IN4(n8277), .IN5(
        n8099), .IN6(n8230), .Q(n8228) );
  NOR2X0 U8252 ( .IN1(n8083), .IN2(n7599), .QN(n7598) );
  AO222X1 U8253 ( .IN1(n8099), .IN2(n8277), .IN3(n8255), .IN4(n7606), .IN5(
        n7609), .IN6(n8256), .Q(n8252) );
  AO222X1 U8254 ( .IN1(n7615), .IN2(n8258), .IN3(n7611), .IN4(n8278), .IN5(
        n7613), .IN6(n8279), .Q(n8256) );
  AO222X1 U8255 ( .IN1(n7613), .IN2(n8278), .IN3(n7615), .IN4(n8257), .IN5(
        n7611), .IN6(n8258), .Q(n8255) );
  AO222X1 U8256 ( .IN1(n7621), .IN2(n8260), .IN3(n7617), .IN4(n8280), .IN5(
        n7619), .IN6(n8281), .Q(n8258) );
  AO222X1 U8257 ( .IN1(n7619), .IN2(n8280), .IN3(n7621), .IN4(n8259), .IN5(
        n7617), .IN6(n8260), .Q(n8257) );
  AO222X1 U8258 ( .IN1(n8262), .IN2(n7626), .IN3(n7623), .IN4(n8282), .IN5(
        n7625), .IN6(n8283), .Q(n8260) );
  AO222X1 U8259 ( .IN1(n7625), .IN2(n8282), .IN3(n8261), .IN4(n7626), .IN5(
        n7623), .IN6(n8262), .Q(n8259) );
  AO222X1 U8260 ( .IN1(n7633), .IN2(n8264), .IN3(n7629), .IN4(n8284), .IN5(
        n7631), .IN6(n8285), .Q(n8262) );
  AO222X1 U8261 ( .IN1(n7631), .IN2(n8284), .IN3(n7633), .IN4(n8263), .IN5(
        n7629), .IN6(n8264), .Q(n8261) );
  AO222X1 U8262 ( .IN1(n8266), .IN2(n7638), .IN3(n7635), .IN4(n8286), .IN5(
        n7637), .IN6(n8287), .Q(n8264) );
  AO222X1 U8263 ( .IN1(n7637), .IN2(n8286), .IN3(n8265), .IN4(n7638), .IN5(
        n7635), .IN6(n8266), .Q(n8263) );
  AO222X1 U8264 ( .IN1(n8268), .IN2(n7644), .IN3(n7641), .IN4(n8288), .IN5(
        n7643), .IN6(n8289), .Q(n8266) );
  AO222X1 U8265 ( .IN1(n7643), .IN2(n8288), .IN3(n8267), .IN4(n7644), .IN5(
        n7641), .IN6(n8268), .Q(n8265) );
  AO222X1 U8266 ( .IN1(n8270), .IN2(n7650), .IN3(n7647), .IN4(n8290), .IN5(
        n7649), .IN6(n8291), .Q(n8268) );
  AO222X1 U8267 ( .IN1(n7649), .IN2(n8290), .IN3(n8269), .IN4(n7650), .IN5(
        n7647), .IN6(n8270), .Q(n8267) );
  AO222X1 U8268 ( .IN1(n7657), .IN2(n8272), .IN3(n7653), .IN4(n8292), .IN5(
        n7655), .IN6(n8293), .Q(n8270) );
  AO222X1 U8269 ( .IN1(n7655), .IN2(n8292), .IN3(n7657), .IN4(n8271), .IN5(
        n7653), .IN6(n8272), .Q(n8269) );
  AO222X1 U8270 ( .IN1(n8274), .IN2(n7660), .IN3(n7659), .IN4(n8294), .IN5(
        n8078), .IN6(n8295), .Q(n8272) );
  AO222X1 U8271 ( .IN1(n8078), .IN2(n8294), .IN3(n8273), .IN4(n7660), .IN5(
        n7659), .IN6(n8274), .Q(n8271) );
  AO222X1 U8272 ( .IN1(n7668), .IN2(n8276), .IN3(n7670), .IN4(n8296), .IN5(
        n8146), .IN6(n8297), .Q(n8274) );
  AO222X1 U8273 ( .IN1(n8146), .IN2(n8296), .IN3(n7668), .IN4(n8275), .IN5(
        n7670), .IN6(n8276), .Q(n8273) );
  AO222X1 U8274 ( .IN1(n7672), .IN2(n7236), .IN3(n7671), .IN4(n7235), .IN5(
        n8225), .IN6(n7237), .Q(n8276) );
  AO222X1 U8275 ( .IN1(n7672), .IN2(n7235), .IN3(n7671), .IN4(n7234), .IN5(
        n8225), .IN6(n7236), .Q(n8275) );
  INVX0 U8276 ( .INP(n3659), .ZN(n7234) );
  INVX0 U8277 ( .INP(n3658), .ZN(n7235) );
  AO222X1 U8278 ( .IN1(n8099), .IN2(n8231), .IN3(n8277), .IN4(n7606), .IN5(
        n7609), .IN6(n8230), .Q(n8229) );
  AO222X1 U8279 ( .IN1(n7615), .IN2(n8279), .IN3(n7611), .IN4(n8298), .IN5(
        n7613), .IN6(n8232), .Q(n8230) );
  NOR2X0 U8280 ( .IN1(n8099), .IN2(n7606), .QN(n7609) );
  AO222X1 U8281 ( .IN1(n7613), .IN2(n8298), .IN3(n7615), .IN4(n8278), .IN5(
        n7611), .IN6(n8279), .Q(n8277) );
  AO222X1 U8282 ( .IN1(n7621), .IN2(n8281), .IN3(n7617), .IN4(n8299), .IN5(
        n7619), .IN6(n8300), .Q(n8279) );
  AO222X1 U8283 ( .IN1(n7619), .IN2(n8299), .IN3(n7621), .IN4(n8280), .IN5(
        n7617), .IN6(n8281), .Q(n8278) );
  AO222X1 U8284 ( .IN1(n8283), .IN2(n7626), .IN3(n7623), .IN4(n8301), .IN5(
        n7625), .IN6(n8302), .Q(n8281) );
  AO222X1 U8285 ( .IN1(n7625), .IN2(n8301), .IN3(n8282), .IN4(n7626), .IN5(
        n7623), .IN6(n8283), .Q(n8280) );
  AO222X1 U8286 ( .IN1(n7633), .IN2(n8285), .IN3(n7629), .IN4(n8303), .IN5(
        n7631), .IN6(n8304), .Q(n8283) );
  AO222X1 U8287 ( .IN1(n7631), .IN2(n8303), .IN3(n7633), .IN4(n8284), .IN5(
        n7629), .IN6(n8285), .Q(n8282) );
  AO222X1 U8288 ( .IN1(n8287), .IN2(n7638), .IN3(n7635), .IN4(n8305), .IN5(
        n7637), .IN6(n8306), .Q(n8285) );
  AO222X1 U8289 ( .IN1(n7637), .IN2(n8305), .IN3(n8286), .IN4(n7638), .IN5(
        n7635), .IN6(n8287), .Q(n8284) );
  AO222X1 U8290 ( .IN1(n8289), .IN2(n7644), .IN3(n7641), .IN4(n8307), .IN5(
        n7643), .IN6(n8308), .Q(n8287) );
  AO222X1 U8291 ( .IN1(n7643), .IN2(n8307), .IN3(n8288), .IN4(n7644), .IN5(
        n7641), .IN6(n8289), .Q(n8286) );
  AO222X1 U8292 ( .IN1(n8291), .IN2(n7650), .IN3(n7647), .IN4(n8309), .IN5(
        n7649), .IN6(n8310), .Q(n8289) );
  AO222X1 U8293 ( .IN1(n7649), .IN2(n8309), .IN3(n8290), .IN4(n7650), .IN5(
        n7647), .IN6(n8291), .Q(n8288) );
  AO222X1 U8294 ( .IN1(n7657), .IN2(n8293), .IN3(n7653), .IN4(n8311), .IN5(
        n7655), .IN6(n8312), .Q(n8291) );
  AO222X1 U8295 ( .IN1(n7655), .IN2(n8311), .IN3(n7657), .IN4(n8292), .IN5(
        n7653), .IN6(n8293), .Q(n8290) );
  AO222X1 U8296 ( .IN1(n8295), .IN2(n7660), .IN3(n7659), .IN4(n8313), .IN5(
        n8078), .IN6(n8314), .Q(n8293) );
  AO222X1 U8297 ( .IN1(n8078), .IN2(n8313), .IN3(n8294), .IN4(n7660), .IN5(
        n7659), .IN6(n8295), .Q(n8292) );
  AO222X1 U8298 ( .IN1(n7668), .IN2(n8297), .IN3(n7670), .IN4(n8315), .IN5(
        n8146), .IN6(n8316), .Q(n8295) );
  AO222X1 U8299 ( .IN1(n8146), .IN2(n8315), .IN3(n7668), .IN4(n8296), .IN5(
        n7670), .IN6(n8297), .Q(n8294) );
  AO222X1 U8300 ( .IN1(n7672), .IN2(n7238), .IN3(n7671), .IN4(n7237), .IN5(
        n8225), .IN6(n7239), .Q(n8297) );
  AO222X1 U8301 ( .IN1(n7672), .IN2(n7237), .IN3(n7671), .IN4(n7236), .IN5(
        n8225), .IN6(n7238), .Q(n8296) );
  INVX0 U8302 ( .INP(n3657), .ZN(n7236) );
  INVX0 U8303 ( .INP(n3656), .ZN(n7237) );
  AO222X1 U8304 ( .IN1(n7613), .IN2(n8233), .IN3(n7615), .IN4(n8298), .IN5(
        n7611), .IN6(n8232), .Q(n8231) );
  AO222X1 U8305 ( .IN1(n7621), .IN2(n8300), .IN3(n7617), .IN4(n8317), .IN5(
        n7619), .IN6(n8234), .Q(n8232) );
  XOR2X1 U8306 ( .IN1(n8318), .IN2(n8319), .Q(n7611) );
  AO222X1 U8307 ( .IN1(n7619), .IN2(n8317), .IN3(n7621), .IN4(n8299), .IN5(
        n7617), .IN6(n8300), .Q(n8298) );
  AO222X1 U8308 ( .IN1(n8302), .IN2(n7626), .IN3(n7623), .IN4(n8320), .IN5(
        n7625), .IN6(n8321), .Q(n8300) );
  AO222X1 U8309 ( .IN1(n7625), .IN2(n8320), .IN3(n8301), .IN4(n7626), .IN5(
        n7623), .IN6(n8302), .Q(n8299) );
  AO222X1 U8310 ( .IN1(n7633), .IN2(n8304), .IN3(n7629), .IN4(n8322), .IN5(
        n7631), .IN6(n8323), .Q(n8302) );
  AO222X1 U8311 ( .IN1(n7631), .IN2(n8322), .IN3(n7633), .IN4(n8303), .IN5(
        n7629), .IN6(n8304), .Q(n8301) );
  AO222X1 U8312 ( .IN1(n8306), .IN2(n7638), .IN3(n7635), .IN4(n8324), .IN5(
        n7637), .IN6(n8325), .Q(n8304) );
  AO222X1 U8313 ( .IN1(n7637), .IN2(n8324), .IN3(n8305), .IN4(n7638), .IN5(
        n7635), .IN6(n8306), .Q(n8303) );
  AO222X1 U8314 ( .IN1(n8308), .IN2(n7644), .IN3(n7641), .IN4(n8326), .IN5(
        n7643), .IN6(n8327), .Q(n8306) );
  AO222X1 U8315 ( .IN1(n7643), .IN2(n8326), .IN3(n8307), .IN4(n7644), .IN5(
        n7641), .IN6(n8308), .Q(n8305) );
  AO222X1 U8316 ( .IN1(n8310), .IN2(n7650), .IN3(n7647), .IN4(n8328), .IN5(
        n7649), .IN6(n8329), .Q(n8308) );
  AO222X1 U8317 ( .IN1(n7649), .IN2(n8328), .IN3(n8309), .IN4(n7650), .IN5(
        n7647), .IN6(n8310), .Q(n8307) );
  AO222X1 U8318 ( .IN1(n7657), .IN2(n8312), .IN3(n7653), .IN4(n8330), .IN5(
        n7655), .IN6(n8331), .Q(n8310) );
  AO222X1 U8319 ( .IN1(n7655), .IN2(n8330), .IN3(n7657), .IN4(n8311), .IN5(
        n7653), .IN6(n8312), .Q(n8309) );
  AO222X1 U8320 ( .IN1(n8314), .IN2(n7660), .IN3(n7659), .IN4(n8332), .IN5(
        n8078), .IN6(n8333), .Q(n8312) );
  AO222X1 U8321 ( .IN1(n8078), .IN2(n8332), .IN3(n8313), .IN4(n7660), .IN5(
        n7659), .IN6(n8314), .Q(n8311) );
  AO222X1 U8322 ( .IN1(n7668), .IN2(n8316), .IN3(n7670), .IN4(n8334), .IN5(
        n8146), .IN6(n8335), .Q(n8314) );
  AO222X1 U8323 ( .IN1(n8146), .IN2(n8334), .IN3(n7668), .IN4(n8315), .IN5(
        n7670), .IN6(n8316), .Q(n8313) );
  AO222X1 U8324 ( .IN1(n7672), .IN2(n7240), .IN3(n7671), .IN4(n7239), .IN5(
        n8225), .IN6(n7241), .Q(n8316) );
  AO222X1 U8325 ( .IN1(n7672), .IN2(n7239), .IN3(n7671), .IN4(n7238), .IN5(
        n8225), .IN6(n7240), .Q(n8315) );
  INVX0 U8326 ( .INP(n3655), .ZN(n7238) );
  INVX0 U8327 ( .INP(n3654), .ZN(n7239) );
  AND2X1 U8328 ( .IN1(n8318), .IN2(n8319), .Q(n7615) );
  AO222X1 U8329 ( .IN1(n7619), .IN2(n8235), .IN3(n7621), .IN4(n8317), .IN5(
        n7617), .IN6(n8234), .Q(n8233) );
  AO222X1 U8330 ( .IN1(n8321), .IN2(n7626), .IN3(n7623), .IN4(n8336), .IN5(
        n7625), .IN6(n8236), .Q(n8234) );
  XOR2X1 U8331 ( .IN1(n8337), .IN2(n8338), .Q(n7617) );
  AO222X1 U8332 ( .IN1(n7625), .IN2(n8336), .IN3(n8320), .IN4(n7626), .IN5(
        n7623), .IN6(n8321), .Q(n8317) );
  AO222X1 U8333 ( .IN1(n7633), .IN2(n8323), .IN3(n7629), .IN4(n8339), .IN5(
        n7631), .IN6(n8340), .Q(n8321) );
  AO222X1 U8334 ( .IN1(n7631), .IN2(n8339), .IN3(n7633), .IN4(n8322), .IN5(
        n7629), .IN6(n8323), .Q(n8320) );
  AO222X1 U8335 ( .IN1(n8325), .IN2(n7638), .IN3(n7635), .IN4(n8341), .IN5(
        n7637), .IN6(n8342), .Q(n8323) );
  AO222X1 U8336 ( .IN1(n7637), .IN2(n8341), .IN3(n8324), .IN4(n7638), .IN5(
        n7635), .IN6(n8325), .Q(n8322) );
  AO222X1 U8337 ( .IN1(n8327), .IN2(n7644), .IN3(n7641), .IN4(n8343), .IN5(
        n7643), .IN6(n8344), .Q(n8325) );
  AO222X1 U8338 ( .IN1(n7643), .IN2(n8343), .IN3(n8326), .IN4(n7644), .IN5(
        n7641), .IN6(n8327), .Q(n8324) );
  AO222X1 U8339 ( .IN1(n8329), .IN2(n7650), .IN3(n7647), .IN4(n8345), .IN5(
        n7649), .IN6(n8346), .Q(n8327) );
  AO222X1 U8340 ( .IN1(n7649), .IN2(n8345), .IN3(n8328), .IN4(n7650), .IN5(
        n7647), .IN6(n8329), .Q(n8326) );
  AO222X1 U8341 ( .IN1(n7657), .IN2(n8331), .IN3(n7653), .IN4(n8347), .IN5(
        n7655), .IN6(n8348), .Q(n8329) );
  AO222X1 U8342 ( .IN1(n7655), .IN2(n8347), .IN3(n7657), .IN4(n8330), .IN5(
        n7653), .IN6(n8331), .Q(n8328) );
  AO222X1 U8343 ( .IN1(n8333), .IN2(n7660), .IN3(n7659), .IN4(n8349), .IN5(
        n8078), .IN6(n8350), .Q(n8331) );
  AO222X1 U8344 ( .IN1(n8078), .IN2(n8349), .IN3(n8332), .IN4(n7660), .IN5(
        n7659), .IN6(n8333), .Q(n8330) );
  AO222X1 U8345 ( .IN1(n7668), .IN2(n8335), .IN3(n7670), .IN4(n8351), .IN5(
        n8146), .IN6(n8352), .Q(n8333) );
  AO222X1 U8346 ( .IN1(n8146), .IN2(n8351), .IN3(n7668), .IN4(n8334), .IN5(
        n7670), .IN6(n8335), .Q(n8332) );
  AO222X1 U8347 ( .IN1(n7672), .IN2(n7242), .IN3(n7671), .IN4(n7241), .IN5(
        n8225), .IN6(n7243), .Q(n8335) );
  AO222X1 U8348 ( .IN1(n7672), .IN2(n7241), .IN3(n7671), .IN4(n7240), .IN5(
        n8225), .IN6(n7242), .Q(n8334) );
  INVX0 U8349 ( .INP(n3653), .ZN(n7240) );
  INVX0 U8350 ( .INP(n3652), .ZN(n7241) );
  NOR2X0 U8351 ( .IN1(n8353), .IN2(n7692), .QN(n7621) );
  AO222X1 U8352 ( .IN1(n7625), .IN2(n8237), .IN3(n8336), .IN4(n7626), .IN5(
        n7623), .IN6(n8236), .Q(n8235) );
  AO222X1 U8353 ( .IN1(n7633), .IN2(n8340), .IN3(n7629), .IN4(n8354), .IN5(
        n7631), .IN6(n8239), .Q(n8236) );
  NOR2X0 U8354 ( .IN1(n7625), .IN2(n7626), .QN(n7623) );
  AO222X1 U8355 ( .IN1(n7631), .IN2(n8354), .IN3(n7633), .IN4(n8339), .IN5(
        n7629), .IN6(n8340), .Q(n8336) );
  AO222X1 U8356 ( .IN1(n8342), .IN2(n7638), .IN3(n7635), .IN4(n8355), .IN5(
        n7637), .IN6(n8356), .Q(n8340) );
  AO222X1 U8357 ( .IN1(n7637), .IN2(n8355), .IN3(n8341), .IN4(n7638), .IN5(
        n7635), .IN6(n8342), .Q(n8339) );
  AO222X1 U8358 ( .IN1(n8344), .IN2(n7644), .IN3(n7641), .IN4(n8357), .IN5(
        n7643), .IN6(n8358), .Q(n8342) );
  AO222X1 U8359 ( .IN1(n7643), .IN2(n8357), .IN3(n8343), .IN4(n7644), .IN5(
        n7641), .IN6(n8344), .Q(n8341) );
  AO222X1 U8360 ( .IN1(n8346), .IN2(n7650), .IN3(n7647), .IN4(n8359), .IN5(
        n7649), .IN6(n8360), .Q(n8344) );
  AO222X1 U8361 ( .IN1(n7649), .IN2(n8359), .IN3(n8345), .IN4(n7650), .IN5(
        n7647), .IN6(n8346), .Q(n8343) );
  AO222X1 U8362 ( .IN1(n7657), .IN2(n8348), .IN3(n7653), .IN4(n8361), .IN5(
        n7655), .IN6(n8362), .Q(n8346) );
  AO222X1 U8363 ( .IN1(n7655), .IN2(n8361), .IN3(n7657), .IN4(n8347), .IN5(
        n7653), .IN6(n8348), .Q(n8345) );
  AO222X1 U8364 ( .IN1(n8350), .IN2(n7660), .IN3(n7659), .IN4(n8363), .IN5(
        n8078), .IN6(n8364), .Q(n8348) );
  AO222X1 U8365 ( .IN1(n8078), .IN2(n8363), .IN3(n8349), .IN4(n7660), .IN5(
        n7659), .IN6(n8350), .Q(n8347) );
  AO222X1 U8366 ( .IN1(n7668), .IN2(n8352), .IN3(n7670), .IN4(n8365), .IN5(
        n8146), .IN6(n8366), .Q(n8350) );
  AO222X1 U8367 ( .IN1(n8146), .IN2(n8365), .IN3(n7668), .IN4(n8351), .IN5(
        n7670), .IN6(n8352), .Q(n8349) );
  AO222X1 U8368 ( .IN1(n7672), .IN2(n7244), .IN3(n7671), .IN4(n7243), .IN5(
        n8225), .IN6(n7245), .Q(n8352) );
  AO222X1 U8369 ( .IN1(n7672), .IN2(n7243), .IN3(n7671), .IN4(n7242), .IN5(
        n8225), .IN6(n7244), .Q(n8351) );
  INVX0 U8370 ( .INP(n3651), .ZN(n7242) );
  INVX0 U8371 ( .INP(n3650), .ZN(n7243) );
  AO222X1 U8372 ( .IN1(n7631), .IN2(n8238), .IN3(n7633), .IN4(n8354), .IN5(
        n7629), .IN6(n8239), .Q(n8237) );
  AO222X1 U8373 ( .IN1(n8356), .IN2(n7638), .IN3(n7635), .IN4(n8367), .IN5(
        n7637), .IN6(n8241), .Q(n8239) );
  XOR2X1 U8374 ( .IN1(n8368), .IN2(n8369), .Q(n7629) );
  AO222X1 U8375 ( .IN1(n7637), .IN2(n8367), .IN3(n8355), .IN4(n7638), .IN5(
        n7635), .IN6(n8356), .Q(n8354) );
  AO222X1 U8376 ( .IN1(n8358), .IN2(n7644), .IN3(n7641), .IN4(n8370), .IN5(
        n7643), .IN6(n8371), .Q(n8356) );
  AO222X1 U8377 ( .IN1(n7643), .IN2(n8370), .IN3(n8357), .IN4(n7644), .IN5(
        n7641), .IN6(n8358), .Q(n8355) );
  AO222X1 U8378 ( .IN1(n8360), .IN2(n7650), .IN3(n7647), .IN4(n8372), .IN5(
        n7649), .IN6(n8373), .Q(n8358) );
  AO222X1 U8379 ( .IN1(n7649), .IN2(n8372), .IN3(n8359), .IN4(n7650), .IN5(
        n7647), .IN6(n8360), .Q(n8357) );
  AO222X1 U8380 ( .IN1(n7657), .IN2(n8362), .IN3(n7653), .IN4(n8374), .IN5(
        n7655), .IN6(n8375), .Q(n8360) );
  AO222X1 U8381 ( .IN1(n7655), .IN2(n8374), .IN3(n7657), .IN4(n8361), .IN5(
        n7653), .IN6(n8362), .Q(n8359) );
  AO222X1 U8382 ( .IN1(n8364), .IN2(n7660), .IN3(n7659), .IN4(n8376), .IN5(
        n8078), .IN6(n8377), .Q(n8362) );
  AO222X1 U8383 ( .IN1(n8078), .IN2(n8376), .IN3(n8363), .IN4(n7660), .IN5(
        n7659), .IN6(n8364), .Q(n8361) );
  AO222X1 U8384 ( .IN1(n7668), .IN2(n8366), .IN3(n7670), .IN4(n8378), .IN5(
        n8146), .IN6(n8379), .Q(n8364) );
  AO222X1 U8385 ( .IN1(n8146), .IN2(n8378), .IN3(n7668), .IN4(n8365), .IN5(
        n7670), .IN6(n8366), .Q(n8363) );
  AO222X1 U8386 ( .IN1(n7672), .IN2(n7246), .IN3(n7671), .IN4(n7245), .IN5(
        n8225), .IN6(n7247), .Q(n8366) );
  AO222X1 U8387 ( .IN1(n7672), .IN2(n7245), .IN3(n7671), .IN4(n7244), .IN5(
        n8225), .IN6(n7246), .Q(n8365) );
  INVX0 U8388 ( .INP(n3649), .ZN(n7244) );
  INVX0 U8389 ( .INP(n3648), .ZN(n7245) );
  NOR2X0 U8390 ( .IN1(n8380), .IN2(n8381), .QN(n7633) );
  AO222X1 U8391 ( .IN1(n8367), .IN2(n7638), .IN3(n7637), .IN4(n8240), .IN5(
        n7635), .IN6(n8241), .Q(n8238) );
  AO222X1 U8392 ( .IN1(n8371), .IN2(n7644), .IN3(n7641), .IN4(n8382), .IN5(
        n7643), .IN6(n8243), .Q(n8241) );
  NOR2X0 U8393 ( .IN1(n7637), .IN2(n7638), .QN(n7635) );
  AO222X1 U8394 ( .IN1(n8382), .IN2(n7644), .IN3(n7643), .IN4(n8242), .IN5(
        n7641), .IN6(n8243), .Q(n8240) );
  AO222X1 U8395 ( .IN1(n8383), .IN2(n7650), .IN3(n7647), .IN4(n8384), .IN5(
        n7649), .IN6(n8245), .Q(n8243) );
  AO222X1 U8396 ( .IN1(n8384), .IN2(n7650), .IN3(n7649), .IN4(n8244), .IN5(
        n7647), .IN6(n8245), .Q(n8242) );
  AO222X1 U8397 ( .IN1(n7657), .IN2(n8385), .IN3(n7653), .IN4(n8386), .IN5(
        n7655), .IN6(n8247), .Q(n8245) );
  AO222X1 U8398 ( .IN1(n7657), .IN2(n8386), .IN3(n7655), .IN4(n8246), .IN5(
        n7653), .IN6(n8247), .Q(n8244) );
  AO222X1 U8399 ( .IN1(n8387), .IN2(n7660), .IN3(n7659), .IN4(n8388), .IN5(
        n8078), .IN6(n8249), .Q(n8247) );
  AO222X1 U8400 ( .IN1(n8388), .IN2(n7660), .IN3(n8078), .IN4(n8248), .IN5(
        n7659), .IN6(n8249), .Q(n8246) );
  AO222X1 U8401 ( .IN1(n7668), .IN2(n8389), .IN3(n7670), .IN4(n8390), .IN5(
        n8146), .IN6(n8251), .Q(n8249) );
  AO222X1 U8402 ( .IN1(n7668), .IN2(n8390), .IN3(n8146), .IN4(n8250), .IN5(
        n7670), .IN6(n8251), .Q(n8248) );
  AO222X1 U8403 ( .IN1(n7672), .IN2(n7258), .IN3(n7671), .IN4(n7257), .IN5(
        n8225), .IN6(n7259), .Q(n8251) );
  AO222X1 U8404 ( .IN1(n7672), .IN2(n7259), .IN3(n7671), .IN4(n7258), .IN5(
        n8225), .IN6(n7260), .Q(n8250) );
  INVX0 U8405 ( .INP(n3633), .ZN(n7260) );
  INVX0 U8406 ( .INP(n3634), .ZN(n7259) );
  INVX0 U8407 ( .INP(n8391), .ZN(n7637) );
  AO222X1 U8408 ( .IN1(n7643), .IN2(n8382), .IN3(n8370), .IN4(n7644), .IN5(
        n7641), .IN6(n8371), .Q(n8367) );
  AO222X1 U8409 ( .IN1(n8373), .IN2(n7650), .IN3(n7647), .IN4(n8392), .IN5(
        n7649), .IN6(n8383), .Q(n8371) );
  NOR2X0 U8410 ( .IN1(n7643), .IN2(n7644), .QN(n7641) );
  AO222X1 U8411 ( .IN1(n7649), .IN2(n8392), .IN3(n8372), .IN4(n7650), .IN5(
        n7647), .IN6(n8373), .Q(n8370) );
  AO222X1 U8412 ( .IN1(n7657), .IN2(n8375), .IN3(n7653), .IN4(n8393), .IN5(
        n7655), .IN6(n8394), .Q(n8373) );
  AO222X1 U8413 ( .IN1(n7655), .IN2(n8393), .IN3(n7657), .IN4(n8374), .IN5(
        n7653), .IN6(n8375), .Q(n8372) );
  AO222X1 U8414 ( .IN1(n8377), .IN2(n7660), .IN3(n7659), .IN4(n8395), .IN5(
        n8078), .IN6(n8396), .Q(n8375) );
  AO222X1 U8415 ( .IN1(n8078), .IN2(n8395), .IN3(n8376), .IN4(n7660), .IN5(
        n7659), .IN6(n8377), .Q(n8374) );
  AO222X1 U8416 ( .IN1(n7668), .IN2(n8379), .IN3(n7670), .IN4(n8397), .IN5(
        n8146), .IN6(n8398), .Q(n8377) );
  AO222X1 U8417 ( .IN1(n8146), .IN2(n8397), .IN3(n7668), .IN4(n8378), .IN5(
        n7670), .IN6(n8379), .Q(n8376) );
  AO222X1 U8418 ( .IN1(n7672), .IN2(n7248), .IN3(n7671), .IN4(n7247), .IN5(
        n8225), .IN6(n7249), .Q(n8379) );
  AO222X1 U8419 ( .IN1(n7672), .IN2(n7247), .IN3(n7671), .IN4(n7246), .IN5(
        n8225), .IN6(n7248), .Q(n8378) );
  INVX0 U8420 ( .INP(n3647), .ZN(n7246) );
  INVX0 U8421 ( .INP(n3646), .ZN(n7247) );
  AO222X1 U8422 ( .IN1(n7649), .IN2(n8384), .IN3(n8392), .IN4(n7650), .IN5(
        n7647), .IN6(n8383), .Q(n8382) );
  AO222X1 U8423 ( .IN1(n7657), .IN2(n8394), .IN3(n7653), .IN4(n8399), .IN5(
        n7655), .IN6(n8385), .Q(n8383) );
  NOR2X0 U8424 ( .IN1(n7649), .IN2(n7650), .QN(n7647) );
  AO222X1 U8425 ( .IN1(n7655), .IN2(n8399), .IN3(n7657), .IN4(n8393), .IN5(
        n7653), .IN6(n8394), .Q(n8392) );
  AO222X1 U8426 ( .IN1(n8396), .IN2(n7660), .IN3(n7659), .IN4(n8400), .IN5(
        n8078), .IN6(n8401), .Q(n8394) );
  AO222X1 U8427 ( .IN1(n8078), .IN2(n8400), .IN3(n8395), .IN4(n7660), .IN5(
        n7659), .IN6(n8396), .Q(n8393) );
  AO222X1 U8428 ( .IN1(n7668), .IN2(n8398), .IN3(n7670), .IN4(n8402), .IN5(
        n8146), .IN6(n8403), .Q(n8396) );
  AO222X1 U8429 ( .IN1(n8146), .IN2(n8402), .IN3(n7668), .IN4(n8397), .IN5(
        n7670), .IN6(n8398), .Q(n8395) );
  AO222X1 U8430 ( .IN1(n7672), .IN2(n7250), .IN3(n7671), .IN4(n7249), .IN5(
        n8225), .IN6(n7251), .Q(n8398) );
  AO222X1 U8431 ( .IN1(n7672), .IN2(n7249), .IN3(n7671), .IN4(n7248), .IN5(
        n8225), .IN6(n7250), .Q(n8397) );
  INVX0 U8432 ( .INP(n3645), .ZN(n7248) );
  INVX0 U8433 ( .INP(n3644), .ZN(n7249) );
  AO222X1 U8434 ( .IN1(n7655), .IN2(n8386), .IN3(n7657), .IN4(n8399), .IN5(
        n7653), .IN6(n8385), .Q(n8384) );
  AO222X1 U8435 ( .IN1(n8401), .IN2(n7660), .IN3(n7659), .IN4(n8404), .IN5(
        n8078), .IN6(n8387), .Q(n8385) );
  XOR2X1 U8436 ( .IN1(n8405), .IN2(n8406), .Q(n7653) );
  AO222X1 U8437 ( .IN1(n8078), .IN2(n8404), .IN3(n8400), .IN4(n7660), .IN5(
        n7659), .IN6(n8401), .Q(n8399) );
  AO222X1 U8438 ( .IN1(n7668), .IN2(n8403), .IN3(n7670), .IN4(n8407), .IN5(
        n8146), .IN6(n8408), .Q(n8401) );
  AO222X1 U8439 ( .IN1(n8146), .IN2(n8407), .IN3(n7668), .IN4(n8402), .IN5(
        n7670), .IN6(n8403), .Q(n8400) );
  AO222X1 U8440 ( .IN1(n7672), .IN2(n7252), .IN3(n7671), .IN4(n7251), .IN5(
        n8225), .IN6(n7253), .Q(n8403) );
  AO222X1 U8441 ( .IN1(n7672), .IN2(n7251), .IN3(n7671), .IN4(n7250), .IN5(
        n8225), .IN6(n7252), .Q(n8402) );
  INVX0 U8442 ( .INP(n3643), .ZN(n7250) );
  INVX0 U8443 ( .INP(n3642), .ZN(n7251) );
  NOR2X0 U8444 ( .IN1(n8409), .IN2(n7681), .QN(n7657) );
  AO222X1 U8445 ( .IN1(n8078), .IN2(n8388), .IN3(n8404), .IN4(n7660), .IN5(
        n7659), .IN6(n8387), .Q(n8386) );
  AO222X1 U8446 ( .IN1(n7668), .IN2(n8408), .IN3(n7670), .IN4(n8410), .IN5(
        n8146), .IN6(n8389), .Q(n8387) );
  NOR2X0 U8447 ( .IN1(n8078), .IN2(n7660), .QN(n7659) );
  AO222X1 U8448 ( .IN1(n8146), .IN2(n8410), .IN3(n7668), .IN4(n8407), .IN5(
        n7670), .IN6(n8408), .Q(n8404) );
  AO222X1 U8449 ( .IN1(n7672), .IN2(n7254), .IN3(n7671), .IN4(n7253), .IN5(
        n8225), .IN6(n7255), .Q(n8408) );
  AO222X1 U8450 ( .IN1(n7672), .IN2(n7253), .IN3(n7671), .IN4(n7252), .IN5(
        n8225), .IN6(n7254), .Q(n8407) );
  INVX0 U8451 ( .INP(n3641), .ZN(n7252) );
  INVX0 U8452 ( .INP(n3640), .ZN(n7253) );
  AO222X1 U8453 ( .IN1(n8146), .IN2(n8390), .IN3(n7668), .IN4(n8410), .IN5(
        n7670), .IN6(n8389), .Q(n8388) );
  AO222X1 U8454 ( .IN1(n7672), .IN2(n7256), .IN3(n7671), .IN4(n7255), .IN5(
        n8225), .IN6(n7257), .Q(n8389) );
  XOR2X1 U8455 ( .IN1(n8411), .IN2(n8412), .Q(n7670) );
  AO222X1 U8456 ( .IN1(n7672), .IN2(n7255), .IN3(n7671), .IN4(n7254), .IN5(
        n8225), .IN6(n7256), .Q(n8410) );
  INVX0 U8457 ( .INP(n3639), .ZN(n7254) );
  INVX0 U8458 ( .INP(n3638), .ZN(n7255) );
  AND2X1 U8459 ( .IN1(n8412), .IN2(n8411), .Q(n7668) );
  AO222X1 U8460 ( .IN1(n7672), .IN2(n7257), .IN3(n7671), .IN4(n7256), .IN5(
        n8225), .IN6(n7258), .Q(n8390) );
  INVX0 U8461 ( .INP(n3635), .ZN(n7258) );
  INVX0 U8462 ( .INP(n3637), .ZN(n7256) );
  INVX0 U8463 ( .INP(n3636), .ZN(n7257) );
  NOR2X0 U8464 ( .IN1(n8225), .IN2(n7671), .QN(n7672) );
  NOR2X0 U8465 ( .IN1(n8411), .IN2(n8412), .QN(n8146) );
  NOR2X0 U8466 ( .IN1(n8405), .IN2(n8406), .QN(n7655) );
  NOR2X0 U8467 ( .IN1(n8368), .IN2(n8369), .QN(n7631) );
  NOR2X0 U8468 ( .IN1(n8338), .IN2(n8337), .QN(n7619) );
  NOR2X0 U8469 ( .IN1(n8319), .IN2(n8318), .QN(n7613) );
  NOR2X0 U8470 ( .IN1(n8254), .IN2(n8253), .QN(n7594) );
  AND2X1 U8471 ( .IN1(n7712), .IN2(n8227), .Q(n7590) );
  OA21X1 U8472 ( .IN1(n8054), .IN2(n8053), .IN3(n7528), .Q(n7581) );
  INVX0 U8473 ( .INP(n8049), .ZN(n7528) );
  NAND3X0 U8474 ( .IN1(n3628), .IN2(n8414), .IN3(n3629), .QN(n8413) );
  NAND2X0 U8475 ( .IN1(n3627), .IN2(n3715), .QN(n8414) );
  INVX0 U8476 ( .INP(n3694), .ZN(n7148) );
  OA21X1 U8477 ( .IN1(n8416), .IN2(n7319), .IN3(n3629), .Q(n8415) );
  INVX0 U8478 ( .INP(n3628), .ZN(n7319) );
  OA21X1 U8479 ( .IN1(n3714), .IN2(n7330), .IN3(n3627), .Q(n8416) );
  INVX0 U8480 ( .INP(n3715), .ZN(n7330) );
  MUX21X1 U8481 ( .IN1(n7298), .IN2(n8417), .S(n8418), .Q(N3015) );
  AO221X1 U8482 ( .IN1(n8419), .IN2(n8417), .IN3(n8418), .IN4(n8420), .IN5(
        n8421), .Q(N3014) );
  AO21X1 U8483 ( .IN1(n8054), .IN2(n7298), .IN3(n8422), .Q(n8421) );
  AO221X1 U8484 ( .IN1(n8419), .IN2(n8420), .IN3(n8418), .IN4(n8423), .IN5(
        n8424), .Q(N3013) );
  AO21X1 U8485 ( .IN1(n8417), .IN2(n8054), .IN3(n8422), .Q(n8424) );
  AO221X1 U8486 ( .IN1(n8419), .IN2(n8423), .IN3(n8418), .IN4(n8425), .IN5(
        n8426), .Q(N3012) );
  AO21X1 U8487 ( .IN1(n8420), .IN2(n8054), .IN3(n8422), .Q(n8426) );
  AO222X1 U8488 ( .IN1(n8427), .IN2(n7684), .IN3(n8417), .IN4(n7683), .IN5(
        n7599), .IN6(n7298), .Q(n8420) );
  AO221X1 U8489 ( .IN1(n8419), .IN2(n8425), .IN3(n8418), .IN4(n8428), .IN5(
        n8429), .Q(N3011) );
  AO21X1 U8490 ( .IN1(n8423), .IN2(n8054), .IN3(n8422), .Q(n8429) );
  AO222X1 U8491 ( .IN1(n7683), .IN2(n8427), .IN3(n8417), .IN4(n7599), .IN5(
        n8430), .IN6(n7684), .Q(n8423) );
  AO221X1 U8492 ( .IN1(n8419), .IN2(n8428), .IN3(n8418), .IN4(n8431), .IN5(
        n8432), .Q(N3010) );
  AO21X1 U8493 ( .IN1(n8425), .IN2(n8054), .IN3(n8422), .Q(n8432) );
  AO222X1 U8494 ( .IN1(n7683), .IN2(n8430), .IN3(n8427), .IN4(n7599), .IN5(
        n8433), .IN6(n7684), .Q(n8425) );
  AO222X1 U8495 ( .IN1(n8434), .IN2(n8435), .IN3(n8417), .IN4(n7690), .IN5(
        n7688), .IN6(n7298), .Q(n8427) );
  AO221X1 U8496 ( .IN1(n8419), .IN2(n8431), .IN3(n8418), .IN4(n8436), .IN5(
        n8437), .Q(N3009) );
  AO21X1 U8497 ( .IN1(n8428), .IN2(n8054), .IN3(n8422), .Q(n8437) );
  AO222X1 U8498 ( .IN1(n7683), .IN2(n8433), .IN3(n8430), .IN4(n7599), .IN5(
        n8438), .IN6(n7684), .Q(n8428) );
  AO222X1 U8499 ( .IN1(n7690), .IN2(n8435), .IN3(n7688), .IN4(n8417), .IN5(
        n8434), .IN6(n8439), .Q(n8430) );
  AO221X1 U8500 ( .IN1(n8419), .IN2(n8436), .IN3(n8418), .IN4(n8440), .IN5(
        n8441), .Q(N3008) );
  AO21X1 U8501 ( .IN1(n8431), .IN2(n8054), .IN3(n8422), .Q(n8441) );
  AO222X1 U8502 ( .IN1(n7683), .IN2(n8438), .IN3(n8433), .IN4(n7599), .IN5(
        n8442), .IN6(n7684), .Q(n8431) );
  AO222X1 U8503 ( .IN1(n7690), .IN2(n8439), .IN3(n7688), .IN4(n8435), .IN5(
        n8434), .IN6(n8443), .Q(n8433) );
  AO221X1 U8504 ( .IN1(n8419), .IN2(n8440), .IN3(n8418), .IN4(n8444), .IN5(
        n8445), .Q(N3007) );
  AO21X1 U8505 ( .IN1(n8436), .IN2(n8054), .IN3(n8422), .Q(n8445) );
  AO222X1 U8506 ( .IN1(n7683), .IN2(n8442), .IN3(n8438), .IN4(n7599), .IN5(
        n8446), .IN6(n7684), .Q(n8436) );
  AO222X1 U8507 ( .IN1(n7690), .IN2(n8443), .IN3(n7688), .IN4(n8439), .IN5(
        n8434), .IN6(n8447), .Q(n8438) );
  AO221X1 U8508 ( .IN1(n8419), .IN2(n8444), .IN3(n8418), .IN4(n8448), .IN5(
        n8449), .Q(N3006) );
  AO21X1 U8509 ( .IN1(n8440), .IN2(n8054), .IN3(n8422), .Q(n8449) );
  AO222X1 U8510 ( .IN1(n7683), .IN2(n8446), .IN3(n8442), .IN4(n7599), .IN5(
        n8450), .IN6(n7684), .Q(n8440) );
  AO222X1 U8511 ( .IN1(n7690), .IN2(n8447), .IN3(n7688), .IN4(n8443), .IN5(
        n8434), .IN6(n8451), .Q(n8442) );
  AO222X1 U8512 ( .IN1(n7698), .IN2(n8439), .IN3(n7694), .IN4(n8435), .IN5(
        n7696), .IN6(n8452), .Q(n8443) );
  AO222X1 U8513 ( .IN1(n7703), .IN2(n8453), .IN3(n8417), .IN4(n7705), .IN5(
        n7701), .IN6(n7298), .Q(n8435) );
  AO221X1 U8514 ( .IN1(n8419), .IN2(n8448), .IN3(n8418), .IN4(n8454), .IN5(
        n8455), .Q(N3005) );
  AO21X1 U8515 ( .IN1(n8444), .IN2(n8054), .IN3(n8422), .Q(n8455) );
  AO222X1 U8516 ( .IN1(n7683), .IN2(n8450), .IN3(n8446), .IN4(n7599), .IN5(
        n8456), .IN6(n7684), .Q(n8444) );
  AO222X1 U8517 ( .IN1(n7690), .IN2(n8451), .IN3(n7688), .IN4(n8447), .IN5(
        n8434), .IN6(n8457), .Q(n8446) );
  AO222X1 U8518 ( .IN1(n7698), .IN2(n8452), .IN3(n7694), .IN4(n8439), .IN5(
        n7696), .IN6(n8458), .Q(n8447) );
  AO222X1 U8519 ( .IN1(n7705), .IN2(n8453), .IN3(n7701), .IN4(n8417), .IN5(
        n7703), .IN6(n8459), .Q(n8439) );
  AO221X1 U8520 ( .IN1(n8419), .IN2(n8454), .IN3(n8418), .IN4(n8460), .IN5(
        n8461), .Q(N3004) );
  AO21X1 U8521 ( .IN1(n8448), .IN2(n8054), .IN3(n8422), .Q(n8461) );
  AO222X1 U8522 ( .IN1(n7683), .IN2(n8456), .IN3(n8450), .IN4(n7599), .IN5(
        n8462), .IN6(n7684), .Q(n8448) );
  AO222X1 U8523 ( .IN1(n7690), .IN2(n8457), .IN3(n7688), .IN4(n8451), .IN5(
        n8434), .IN6(n8463), .Q(n8450) );
  AO222X1 U8524 ( .IN1(n7698), .IN2(n8458), .IN3(n7694), .IN4(n8452), .IN5(
        n7696), .IN6(n8464), .Q(n8451) );
  AO222X1 U8525 ( .IN1(n7705), .IN2(n8459), .IN3(n7701), .IN4(n8453), .IN5(
        n7703), .IN6(n8465), .Q(n8452) );
  AO222X1 U8526 ( .IN1(n7716), .IN2(n8466), .IN3(n8417), .IN4(n7714), .IN5(
        n7718), .IN6(n7298), .Q(n8453) );
  AO221X1 U8527 ( .IN1(n8419), .IN2(n8460), .IN3(n8418), .IN4(n8467), .IN5(
        n8468), .Q(N3003) );
  AO21X1 U8528 ( .IN1(n8454), .IN2(n8054), .IN3(n8422), .Q(n8468) );
  AO222X1 U8529 ( .IN1(n7683), .IN2(n8462), .IN3(n8456), .IN4(n7599), .IN5(
        n8469), .IN6(n7684), .Q(n8454) );
  AO222X1 U8530 ( .IN1(n7690), .IN2(n8463), .IN3(n7688), .IN4(n8457), .IN5(
        n8434), .IN6(n8470), .Q(n8456) );
  AO222X1 U8531 ( .IN1(n7698), .IN2(n8464), .IN3(n7694), .IN4(n8458), .IN5(
        n7696), .IN6(n8471), .Q(n8457) );
  AO222X1 U8532 ( .IN1(n7705), .IN2(n8465), .IN3(n7701), .IN4(n8459), .IN5(
        n7703), .IN6(n8472), .Q(n8458) );
  AO222X1 U8533 ( .IN1(n7714), .IN2(n8466), .IN3(n7718), .IN4(n8417), .IN5(
        n7716), .IN6(n8473), .Q(n8459) );
  MUX21X1 U8534 ( .IN1(n7298), .IN2(n8474), .S(n7745), .Q(n8417) );
  AO221X1 U8535 ( .IN1(n8419), .IN2(n8467), .IN3(n8418), .IN4(n8475), .IN5(
        n8476), .Q(N3002) );
  AO21X1 U8536 ( .IN1(n8460), .IN2(n8054), .IN3(n8422), .Q(n8476) );
  AO222X1 U8537 ( .IN1(n7683), .IN2(n8469), .IN3(n8462), .IN4(n7599), .IN5(
        n8477), .IN6(n7684), .Q(n8460) );
  AO222X1 U8538 ( .IN1(n7690), .IN2(n8470), .IN3(n7688), .IN4(n8463), .IN5(
        n8434), .IN6(n8478), .Q(n8462) );
  AO222X1 U8539 ( .IN1(n7698), .IN2(n8471), .IN3(n7694), .IN4(n8464), .IN5(
        n7696), .IN6(n8479), .Q(n8463) );
  AO222X1 U8540 ( .IN1(n7705), .IN2(n8472), .IN3(n7701), .IN4(n8465), .IN5(
        n7703), .IN6(n8480), .Q(n8464) );
  AO222X1 U8541 ( .IN1(n7714), .IN2(n8473), .IN3(n7718), .IN4(n8466), .IN5(
        n7716), .IN6(n8481), .Q(n8465) );
  AO221X1 U8542 ( .IN1(n8419), .IN2(n8475), .IN3(n8418), .IN4(n8482), .IN5(
        n8483), .Q(N3001) );
  AO21X1 U8543 ( .IN1(n8467), .IN2(n8054), .IN3(n8422), .Q(n8483) );
  AO222X1 U8544 ( .IN1(n7683), .IN2(n8477), .IN3(n8469), .IN4(n7599), .IN5(
        n8484), .IN6(n7684), .Q(n8467) );
  AO222X1 U8545 ( .IN1(n7690), .IN2(n8478), .IN3(n7688), .IN4(n8470), .IN5(
        n8434), .IN6(n8485), .Q(n8469) );
  AO222X1 U8546 ( .IN1(n7698), .IN2(n8479), .IN3(n7694), .IN4(n8471), .IN5(
        n7696), .IN6(n8486), .Q(n8470) );
  AO222X1 U8547 ( .IN1(n7705), .IN2(n8480), .IN3(n7701), .IN4(n8472), .IN5(
        n7703), .IN6(n8487), .Q(n8471) );
  AO221X1 U8548 ( .IN1(n8419), .IN2(n8482), .IN3(n8418), .IN4(n8488), .IN5(
        n8489), .Q(N3000) );
  AO21X1 U8549 ( .IN1(n8475), .IN2(n8054), .IN3(n8422), .Q(n8489) );
  AO222X1 U8550 ( .IN1(n7683), .IN2(n8484), .IN3(n8477), .IN4(n7599), .IN5(
        n8490), .IN6(n7684), .Q(n8475) );
  AO222X1 U8551 ( .IN1(n7690), .IN2(n8485), .IN3(n7688), .IN4(n8478), .IN5(
        n8434), .IN6(n8491), .Q(n8477) );
  AO222X1 U8552 ( .IN1(n7698), .IN2(n8486), .IN3(n7694), .IN4(n8479), .IN5(
        n7696), .IN6(n8492), .Q(n8478) );
  AO222X1 U8553 ( .IN1(n7705), .IN2(n8487), .IN3(n7701), .IN4(n8480), .IN5(
        n7703), .IN6(n8493), .Q(n8479) );
  AO221X1 U8554 ( .IN1(n8419), .IN2(n8488), .IN3(n8418), .IN4(n8494), .IN5(
        n8495), .Q(N2999) );
  AO21X1 U8555 ( .IN1(n8482), .IN2(n8054), .IN3(n8422), .Q(n8495) );
  AO222X1 U8556 ( .IN1(n7683), .IN2(n8490), .IN3(n8484), .IN4(n7599), .IN5(
        n8496), .IN6(n7684), .Q(n8482) );
  AO222X1 U8557 ( .IN1(n7690), .IN2(n8491), .IN3(n7688), .IN4(n8485), .IN5(
        n8434), .IN6(n8497), .Q(n8484) );
  AO222X1 U8558 ( .IN1(n7698), .IN2(n8492), .IN3(n7694), .IN4(n8486), .IN5(
        n7696), .IN6(n8498), .Q(n8485) );
  AO222X1 U8559 ( .IN1(n7705), .IN2(n8493), .IN3(n7701), .IN4(n8487), .IN5(
        n7703), .IN6(n8499), .Q(n8486) );
  AO222X1 U8560 ( .IN1(n8500), .IN2(n8480), .IN3(n7709), .IN4(n8472), .IN5(
        n8501), .IN6(n8502), .Q(n8487) );
  AO222X1 U8561 ( .IN1(n7714), .IN2(n8481), .IN3(n7718), .IN4(n8473), .IN5(
        n7716), .IN6(n8503), .Q(n8472) );
  AO221X1 U8562 ( .IN1(n8419), .IN2(n8494), .IN3(n8418), .IN4(n8504), .IN5(
        n8505), .Q(N2998) );
  AO21X1 U8563 ( .IN1(n8488), .IN2(n8054), .IN3(n8422), .Q(n8505) );
  AO222X1 U8564 ( .IN1(n7683), .IN2(n8496), .IN3(n8490), .IN4(n7599), .IN5(
        n8506), .IN6(n7684), .Q(n8488) );
  AO222X1 U8565 ( .IN1(n7690), .IN2(n8497), .IN3(n7688), .IN4(n8491), .IN5(
        n8434), .IN6(n8507), .Q(n8490) );
  AO222X1 U8566 ( .IN1(n7698), .IN2(n8498), .IN3(n7694), .IN4(n8492), .IN5(
        n7696), .IN6(n8508), .Q(n8491) );
  AO222X1 U8567 ( .IN1(n7705), .IN2(n8499), .IN3(n7701), .IN4(n8493), .IN5(
        n7703), .IN6(n8509), .Q(n8492) );
  AO222X1 U8568 ( .IN1(n8500), .IN2(n8502), .IN3(n7709), .IN4(n8480), .IN5(
        n8501), .IN6(n8510), .Q(n8493) );
  AO222X1 U8569 ( .IN1(n7714), .IN2(n8503), .IN3(n7718), .IN4(n8481), .IN5(
        n7716), .IN6(n8511), .Q(n8480) );
  AO222X1 U8570 ( .IN1(n7720), .IN2(n8473), .IN3(n7724), .IN4(n8466), .IN5(
        n7722), .IN6(n8512), .Q(n8481) );
  AO222X1 U8571 ( .IN1(n7745), .IN2(n8513), .IN3(n8474), .IN4(n7743), .IN5(
        n7747), .IN6(n7298), .Q(n8466) );
  AO221X1 U8572 ( .IN1(n8419), .IN2(n8504), .IN3(n8418), .IN4(n8514), .IN5(
        n8515), .Q(N2997) );
  AO21X1 U8573 ( .IN1(n8494), .IN2(n8054), .IN3(n8422), .Q(n8515) );
  AO222X1 U8574 ( .IN1(n7683), .IN2(n8506), .IN3(n8496), .IN4(n7599), .IN5(
        n8516), .IN6(n7684), .Q(n8494) );
  AO222X1 U8575 ( .IN1(n7690), .IN2(n8507), .IN3(n7688), .IN4(n8497), .IN5(
        n8434), .IN6(n8517), .Q(n8496) );
  AO222X1 U8576 ( .IN1(n7698), .IN2(n8508), .IN3(n7694), .IN4(n8498), .IN5(
        n7696), .IN6(n8518), .Q(n8497) );
  AO222X1 U8577 ( .IN1(n7705), .IN2(n8509), .IN3(n7701), .IN4(n8499), .IN5(
        n7703), .IN6(n8519), .Q(n8498) );
  AO222X1 U8578 ( .IN1(n8500), .IN2(n8510), .IN3(n7709), .IN4(n8502), .IN5(
        n8501), .IN6(n8520), .Q(n8499) );
  AO222X1 U8579 ( .IN1(n7714), .IN2(n8511), .IN3(n7718), .IN4(n8503), .IN5(
        n7716), .IN6(n8521), .Q(n8502) );
  AO222X1 U8580 ( .IN1(n7720), .IN2(n8512), .IN3(n7724), .IN4(n8473), .IN5(
        n7722), .IN6(n8522), .Q(n8503) );
  AO222X1 U8581 ( .IN1(n7743), .IN2(n8513), .IN3(n7747), .IN4(n8474), .IN5(
        n7745), .IN6(n8523), .Q(n8473) );
  MUX21X1 U8582 ( .IN1(n7298), .IN2(n8524), .S(n8525), .Q(n8474) );
  AO221X1 U8583 ( .IN1(n8419), .IN2(n8514), .IN3(n8418), .IN4(n8526), .IN5(
        n8527), .Q(N2996) );
  AO21X1 U8584 ( .IN1(n8504), .IN2(n8054), .IN3(n8422), .Q(n8527) );
  AO222X1 U8585 ( .IN1(n7683), .IN2(n8516), .IN3(n8506), .IN4(n7599), .IN5(
        n8528), .IN6(n7684), .Q(n8504) );
  AO222X1 U8586 ( .IN1(n7690), .IN2(n8517), .IN3(n7688), .IN4(n8507), .IN5(
        n8434), .IN6(n8529), .Q(n8506) );
  AO222X1 U8587 ( .IN1(n7698), .IN2(n8518), .IN3(n7694), .IN4(n8508), .IN5(
        n7696), .IN6(n8530), .Q(n8507) );
  AO222X1 U8588 ( .IN1(n7705), .IN2(n8519), .IN3(n7701), .IN4(n8509), .IN5(
        n7703), .IN6(n8531), .Q(n8508) );
  AO222X1 U8589 ( .IN1(n8500), .IN2(n8520), .IN3(n7709), .IN4(n8510), .IN5(
        n8501), .IN6(n8532), .Q(n8509) );
  AO222X1 U8590 ( .IN1(n7714), .IN2(n8521), .IN3(n7718), .IN4(n8511), .IN5(
        n7716), .IN6(n8533), .Q(n8510) );
  AO222X1 U8591 ( .IN1(n7720), .IN2(n8522), .IN3(n7724), .IN4(n8512), .IN5(
        n7722), .IN6(n8534), .Q(n8511) );
  AO222X1 U8592 ( .IN1(n7743), .IN2(n8523), .IN3(n7747), .IN4(n8513), .IN5(
        n7745), .IN6(n8535), .Q(n8512) );
  AO222X1 U8593 ( .IN1(n8524), .IN2(n8536), .IN3(n8525), .IN4(n8537), .IN5(
        n8538), .IN6(n7298), .Q(n8513) );
  AO221X1 U8594 ( .IN1(n8419), .IN2(n8526), .IN3(n8418), .IN4(n8539), .IN5(
        n8540), .Q(N2995) );
  AO21X1 U8595 ( .IN1(n8514), .IN2(n8054), .IN3(n8422), .Q(n8540) );
  AO222X1 U8596 ( .IN1(n7683), .IN2(n8528), .IN3(n8516), .IN4(n7599), .IN5(
        n8541), .IN6(n7684), .Q(n8514) );
  AO222X1 U8597 ( .IN1(n7690), .IN2(n8529), .IN3(n7688), .IN4(n8517), .IN5(
        n8434), .IN6(n8542), .Q(n8516) );
  AO222X1 U8598 ( .IN1(n7698), .IN2(n8530), .IN3(n7694), .IN4(n8518), .IN5(
        n7696), .IN6(n8543), .Q(n8517) );
  AO222X1 U8599 ( .IN1(n7705), .IN2(n8531), .IN3(n7701), .IN4(n8519), .IN5(
        n7703), .IN6(n8544), .Q(n8518) );
  AO222X1 U8600 ( .IN1(n8500), .IN2(n8532), .IN3(n7709), .IN4(n8520), .IN5(
        n8501), .IN6(n8545), .Q(n8519) );
  AO222X1 U8601 ( .IN1(n7714), .IN2(n8533), .IN3(n7718), .IN4(n8521), .IN5(
        n7716), .IN6(n8546), .Q(n8520) );
  AO222X1 U8602 ( .IN1(n7720), .IN2(n8534), .IN3(n7724), .IN4(n8522), .IN5(
        n7722), .IN6(n8547), .Q(n8521) );
  AO221X1 U8603 ( .IN1(n8419), .IN2(n8539), .IN3(n8418), .IN4(n8548), .IN5(
        n8549), .Q(N2994) );
  AO21X1 U8604 ( .IN1(n8526), .IN2(n8054), .IN3(n8422), .Q(n8549) );
  AO222X1 U8605 ( .IN1(n7683), .IN2(n8541), .IN3(n8528), .IN4(n7599), .IN5(
        n8550), .IN6(n7684), .Q(n8526) );
  AO222X1 U8606 ( .IN1(n7690), .IN2(n8542), .IN3(n7688), .IN4(n8529), .IN5(
        n8434), .IN6(n8551), .Q(n8528) );
  AO222X1 U8607 ( .IN1(n7698), .IN2(n8543), .IN3(n7694), .IN4(n8530), .IN5(
        n7696), .IN6(n8552), .Q(n8529) );
  AO222X1 U8608 ( .IN1(n7705), .IN2(n8544), .IN3(n7701), .IN4(n8531), .IN5(
        n7703), .IN6(n8553), .Q(n8530) );
  AO222X1 U8609 ( .IN1(n8500), .IN2(n8545), .IN3(n7709), .IN4(n8532), .IN5(
        n8501), .IN6(n8554), .Q(n8531) );
  AO222X1 U8610 ( .IN1(n7714), .IN2(n8546), .IN3(n7718), .IN4(n8533), .IN5(
        n7716), .IN6(n8555), .Q(n8532) );
  AO222X1 U8611 ( .IN1(n7720), .IN2(n8547), .IN3(n7724), .IN4(n8534), .IN5(
        n7722), .IN6(n8556), .Q(n8533) );
  AO221X1 U8612 ( .IN1(n8419), .IN2(n8548), .IN3(n8418), .IN4(n8557), .IN5(
        n8558), .Q(N2993) );
  AO21X1 U8613 ( .IN1(n8539), .IN2(n8054), .IN3(n8422), .Q(n8558) );
  AO222X1 U8614 ( .IN1(n7683), .IN2(n8550), .IN3(n8541), .IN4(n7599), .IN5(
        n8559), .IN6(n7684), .Q(n8539) );
  AO222X1 U8615 ( .IN1(n7690), .IN2(n8551), .IN3(n7688), .IN4(n8542), .IN5(
        n8434), .IN6(n8560), .Q(n8541) );
  AO222X1 U8616 ( .IN1(n7698), .IN2(n8552), .IN3(n7694), .IN4(n8543), .IN5(
        n7696), .IN6(n8561), .Q(n8542) );
  AO222X1 U8617 ( .IN1(n7705), .IN2(n8553), .IN3(n7701), .IN4(n8544), .IN5(
        n7703), .IN6(n8562), .Q(n8543) );
  AO222X1 U8618 ( .IN1(n8500), .IN2(n8554), .IN3(n7709), .IN4(n8545), .IN5(
        n8501), .IN6(n8563), .Q(n8544) );
  AO222X1 U8619 ( .IN1(n7714), .IN2(n8555), .IN3(n7718), .IN4(n8546), .IN5(
        n7716), .IN6(n8564), .Q(n8545) );
  AO222X1 U8620 ( .IN1(n7720), .IN2(n8556), .IN3(n7724), .IN4(n8547), .IN5(
        n7722), .IN6(n8565), .Q(n8546) );
  AO222X1 U8621 ( .IN1(n7728), .IN2(n8534), .IN3(n7733), .IN4(n8522), .IN5(
        n8566), .IN6(n8567), .Q(n8547) );
  AO222X1 U8622 ( .IN1(n7743), .IN2(n8535), .IN3(n7747), .IN4(n8523), .IN5(
        n7745), .IN6(n8568), .Q(n8522) );
  AO221X1 U8623 ( .IN1(n8419), .IN2(n8557), .IN3(n8418), .IN4(n8569), .IN5(
        n8570), .Q(N2992) );
  AO21X1 U8624 ( .IN1(n8548), .IN2(n8054), .IN3(n8422), .Q(n8570) );
  AO222X1 U8625 ( .IN1(n7683), .IN2(n8559), .IN3(n8550), .IN4(n7599), .IN5(
        n8571), .IN6(n7684), .Q(n8548) );
  AO222X1 U8626 ( .IN1(n7690), .IN2(n8560), .IN3(n7688), .IN4(n8551), .IN5(
        n8434), .IN6(n8572), .Q(n8550) );
  AO222X1 U8627 ( .IN1(n7698), .IN2(n8561), .IN3(n7694), .IN4(n8552), .IN5(
        n7696), .IN6(n8573), .Q(n8551) );
  AO222X1 U8628 ( .IN1(n7705), .IN2(n8562), .IN3(n7701), .IN4(n8553), .IN5(
        n7703), .IN6(n8574), .Q(n8552) );
  AO222X1 U8629 ( .IN1(n8500), .IN2(n8563), .IN3(n7709), .IN4(n8554), .IN5(
        n8501), .IN6(n8575), .Q(n8553) );
  AO222X1 U8630 ( .IN1(n7714), .IN2(n8564), .IN3(n7718), .IN4(n8555), .IN5(
        n7716), .IN6(n8576), .Q(n8554) );
  AO222X1 U8631 ( .IN1(n7720), .IN2(n8565), .IN3(n7724), .IN4(n8556), .IN5(
        n7722), .IN6(n8577), .Q(n8555) );
  AO222X1 U8632 ( .IN1(n7728), .IN2(n8567), .IN3(n7733), .IN4(n8534), .IN5(
        n8566), .IN6(n8578), .Q(n8556) );
  AO221X1 U8633 ( .IN1(n8419), .IN2(n8569), .IN3(n8418), .IN4(n8579), .IN5(
        n8580), .Q(N2991) );
  AO21X1 U8634 ( .IN1(n8557), .IN2(n8054), .IN3(n8422), .Q(n8580) );
  AO222X1 U8635 ( .IN1(n7683), .IN2(n8571), .IN3(n8559), .IN4(n7599), .IN5(
        n8581), .IN6(n7684), .Q(n8557) );
  AO222X1 U8636 ( .IN1(n7690), .IN2(n8572), .IN3(n7688), .IN4(n8560), .IN5(
        n8434), .IN6(n8582), .Q(n8559) );
  AO222X1 U8637 ( .IN1(n7698), .IN2(n8573), .IN3(n7694), .IN4(n8561), .IN5(
        n7696), .IN6(n8583), .Q(n8560) );
  AO222X1 U8638 ( .IN1(n7705), .IN2(n8574), .IN3(n7701), .IN4(n8562), .IN5(
        n7703), .IN6(n8584), .Q(n8561) );
  AO222X1 U8639 ( .IN1(n8500), .IN2(n8575), .IN3(n7709), .IN4(n8563), .IN5(
        n8501), .IN6(n8585), .Q(n8562) );
  AO222X1 U8640 ( .IN1(n7714), .IN2(n8576), .IN3(n7718), .IN4(n8564), .IN5(
        n7716), .IN6(n8586), .Q(n8563) );
  AO222X1 U8641 ( .IN1(n7720), .IN2(n8577), .IN3(n7724), .IN4(n8565), .IN5(
        n7722), .IN6(n8587), .Q(n8564) );
  AO222X1 U8642 ( .IN1(n7728), .IN2(n8578), .IN3(n7733), .IN4(n8567), .IN5(
        n8566), .IN6(n8588), .Q(n8565) );
  AO221X1 U8643 ( .IN1(n8419), .IN2(n8579), .IN3(n8418), .IN4(n8589), .IN5(
        n8590), .Q(N2990) );
  AO21X1 U8644 ( .IN1(n8569), .IN2(n8054), .IN3(n8422), .Q(n8590) );
  AO222X1 U8645 ( .IN1(n7683), .IN2(n8581), .IN3(n8571), .IN4(n7599), .IN5(
        n8591), .IN6(n7684), .Q(n8569) );
  AO222X1 U8646 ( .IN1(n7690), .IN2(n8582), .IN3(n7688), .IN4(n8572), .IN5(
        n8434), .IN6(n8592), .Q(n8571) );
  AO222X1 U8647 ( .IN1(n7698), .IN2(n8583), .IN3(n7694), .IN4(n8573), .IN5(
        n7696), .IN6(n8593), .Q(n8572) );
  AO222X1 U8648 ( .IN1(n7705), .IN2(n8584), .IN3(n7701), .IN4(n8574), .IN5(
        n7703), .IN6(n8594), .Q(n8573) );
  AO222X1 U8649 ( .IN1(n8500), .IN2(n8585), .IN3(n7709), .IN4(n8575), .IN5(
        n8501), .IN6(n8595), .Q(n8574) );
  AO222X1 U8650 ( .IN1(n7714), .IN2(n8586), .IN3(n7718), .IN4(n8576), .IN5(
        n7716), .IN6(n8596), .Q(n8575) );
  AO222X1 U8651 ( .IN1(n7720), .IN2(n8587), .IN3(n7724), .IN4(n8577), .IN5(
        n7722), .IN6(n8597), .Q(n8576) );
  AO222X1 U8652 ( .IN1(n7728), .IN2(n8588), .IN3(n7733), .IN4(n8578), .IN5(
        n8566), .IN6(n8598), .Q(n8577) );
  AO222X1 U8653 ( .IN1(n7737), .IN2(n8567), .IN3(n7741), .IN4(n8534), .IN5(
        n7739), .IN6(n8599), .Q(n8578) );
  AO222X1 U8654 ( .IN1(n7743), .IN2(n8568), .IN3(n7747), .IN4(n8535), .IN5(
        n7745), .IN6(n8600), .Q(n8534) );
  AO221X1 U8655 ( .IN1(n8419), .IN2(n8589), .IN3(n8418), .IN4(n8601), .IN5(
        n8602), .Q(N2989) );
  AO21X1 U8656 ( .IN1(n8579), .IN2(n8054), .IN3(n8422), .Q(n8602) );
  AO222X1 U8657 ( .IN1(n7683), .IN2(n8591), .IN3(n8581), .IN4(n7599), .IN5(
        n8603), .IN6(n7684), .Q(n8579) );
  AO222X1 U8658 ( .IN1(n7690), .IN2(n8592), .IN3(n7688), .IN4(n8582), .IN5(
        n8434), .IN6(n8604), .Q(n8581) );
  AO222X1 U8659 ( .IN1(n7698), .IN2(n8593), .IN3(n7694), .IN4(n8583), .IN5(
        n7696), .IN6(n8605), .Q(n8582) );
  AO222X1 U8660 ( .IN1(n7705), .IN2(n8594), .IN3(n7701), .IN4(n8584), .IN5(
        n7703), .IN6(n8606), .Q(n8583) );
  AO222X1 U8661 ( .IN1(n8500), .IN2(n8595), .IN3(n7709), .IN4(n8585), .IN5(
        n8501), .IN6(n8607), .Q(n8584) );
  AO222X1 U8662 ( .IN1(n7714), .IN2(n8596), .IN3(n7718), .IN4(n8586), .IN5(
        n7716), .IN6(n8608), .Q(n8585) );
  AO222X1 U8663 ( .IN1(n7720), .IN2(n8597), .IN3(n7724), .IN4(n8587), .IN5(
        n7722), .IN6(n8609), .Q(n8586) );
  AO222X1 U8664 ( .IN1(n7728), .IN2(n8598), .IN3(n7733), .IN4(n8588), .IN5(
        n8566), .IN6(n8610), .Q(n8587) );
  AO222X1 U8665 ( .IN1(n7737), .IN2(n8599), .IN3(n7741), .IN4(n8567), .IN5(
        n7739), .IN6(n8611), .Q(n8588) );
  AO222X1 U8666 ( .IN1(n7743), .IN2(n8600), .IN3(n7747), .IN4(n8568), .IN5(
        n7745), .IN6(n8612), .Q(n8567) );
  AO221X1 U8667 ( .IN1(n8419), .IN2(n8601), .IN3(n8418), .IN4(n8613), .IN5(
        n8614), .Q(N2988) );
  AO21X1 U8668 ( .IN1(n8589), .IN2(n8054), .IN3(n8422), .Q(n8614) );
  AO222X1 U8669 ( .IN1(n7683), .IN2(n8603), .IN3(n8591), .IN4(n7599), .IN5(
        n8615), .IN6(n7684), .Q(n8589) );
  AO222X1 U8670 ( .IN1(n7690), .IN2(n8604), .IN3(n7688), .IN4(n8592), .IN5(
        n8434), .IN6(n8616), .Q(n8591) );
  AO222X1 U8671 ( .IN1(n7698), .IN2(n8605), .IN3(n7694), .IN4(n8593), .IN5(
        n7696), .IN6(n8617), .Q(n8592) );
  AO222X1 U8672 ( .IN1(n7705), .IN2(n8606), .IN3(n7701), .IN4(n8594), .IN5(
        n7703), .IN6(n8618), .Q(n8593) );
  AO222X1 U8673 ( .IN1(n8500), .IN2(n8607), .IN3(n7709), .IN4(n8595), .IN5(
        n8501), .IN6(n8619), .Q(n8594) );
  AO222X1 U8674 ( .IN1(n7714), .IN2(n8608), .IN3(n7718), .IN4(n8596), .IN5(
        n7716), .IN6(n8620), .Q(n8595) );
  AO222X1 U8675 ( .IN1(n7720), .IN2(n8609), .IN3(n7724), .IN4(n8597), .IN5(
        n7722), .IN6(n8621), .Q(n8596) );
  AO222X1 U8676 ( .IN1(n7728), .IN2(n8610), .IN3(n7733), .IN4(n8598), .IN5(
        n8566), .IN6(n8622), .Q(n8597) );
  AO221X1 U8677 ( .IN1(n8419), .IN2(n8613), .IN3(n8418), .IN4(n8623), .IN5(
        n8624), .Q(N2987) );
  AO21X1 U8678 ( .IN1(n8601), .IN2(n8054), .IN3(n8422), .Q(n8624) );
  AO222X1 U8679 ( .IN1(n7683), .IN2(n8615), .IN3(n8603), .IN4(n7599), .IN5(
        n8625), .IN6(n7684), .Q(n8601) );
  AO222X1 U8680 ( .IN1(n7690), .IN2(n8616), .IN3(n7688), .IN4(n8604), .IN5(
        n8434), .IN6(n8626), .Q(n8603) );
  AO222X1 U8681 ( .IN1(n7698), .IN2(n8617), .IN3(n7694), .IN4(n8605), .IN5(
        n7696), .IN6(n8627), .Q(n8604) );
  AO222X1 U8682 ( .IN1(n7705), .IN2(n8618), .IN3(n7701), .IN4(n8606), .IN5(
        n7703), .IN6(n8628), .Q(n8605) );
  AO222X1 U8683 ( .IN1(n8500), .IN2(n8619), .IN3(n7709), .IN4(n8607), .IN5(
        n8501), .IN6(n8629), .Q(n8606) );
  AO222X1 U8684 ( .IN1(n7714), .IN2(n8620), .IN3(n7718), .IN4(n8608), .IN5(
        n7716), .IN6(n8630), .Q(n8607) );
  AO222X1 U8685 ( .IN1(n7720), .IN2(n8621), .IN3(n7724), .IN4(n8609), .IN5(
        n7722), .IN6(n8631), .Q(n8608) );
  AO222X1 U8686 ( .IN1(n7728), .IN2(n8622), .IN3(n7733), .IN4(n8610), .IN5(
        n8566), .IN6(n8632), .Q(n8609) );
  AO221X1 U8687 ( .IN1(n8418), .IN2(n8633), .IN3(n8419), .IN4(n8623), .IN5(
        n8634), .Q(N2986) );
  AO21X1 U8688 ( .IN1(n8613), .IN2(n8054), .IN3(n8422), .Q(n8634) );
  AO222X1 U8689 ( .IN1(n8635), .IN2(n7684), .IN3(n8615), .IN4(n7599), .IN5(
        n7683), .IN6(n8625), .Q(n8613) );
  AO222X1 U8690 ( .IN1(n8434), .IN2(n8636), .IN3(n7688), .IN4(n8616), .IN5(
        n7690), .IN6(n8626), .Q(n8615) );
  AO222X1 U8691 ( .IN1(n7696), .IN2(n8637), .IN3(n7694), .IN4(n8617), .IN5(
        n7698), .IN6(n8627), .Q(n8616) );
  AO222X1 U8692 ( .IN1(n7703), .IN2(n8638), .IN3(n7701), .IN4(n8618), .IN5(
        n7705), .IN6(n8628), .Q(n8617) );
  AO222X1 U8693 ( .IN1(n8501), .IN2(n8639), .IN3(n7709), .IN4(n8619), .IN5(
        n8500), .IN6(n8629), .Q(n8618) );
  AO222X1 U8694 ( .IN1(n7716), .IN2(n8640), .IN3(n7718), .IN4(n8620), .IN5(
        n7714), .IN6(n8630), .Q(n8619) );
  AO222X1 U8695 ( .IN1(n7722), .IN2(n8641), .IN3(n7724), .IN4(n8621), .IN5(
        n7720), .IN6(n8631), .Q(n8620) );
  AO222X1 U8696 ( .IN1(n8566), .IN2(n8642), .IN3(n7733), .IN4(n8622), .IN5(
        n7728), .IN6(n8632), .Q(n8621) );
  AO222X1 U8697 ( .IN1(n8099), .IN2(n8643), .IN3(n8598), .IN4(n8254), .IN5(
        n7730), .IN6(n8610), .Q(n8622) );
  AO222X1 U8698 ( .IN1(n7739), .IN2(n8644), .IN3(n7741), .IN4(n8599), .IN5(
        n7737), .IN6(n8611), .Q(n8598) );
  AO222X1 U8699 ( .IN1(n7745), .IN2(n8645), .IN3(n7747), .IN4(n8600), .IN5(
        n7743), .IN6(n8612), .Q(n8599) );
  AO222X1 U8700 ( .IN1(n7643), .IN2(n8646), .IN3(n8535), .IN4(n7626), .IN5(
        n8647), .IN6(n8568), .Q(n8600) );
  AO221X1 U8701 ( .IN1(n8623), .IN2(n8054), .IN3(n8418), .IN4(n7691), .IN5(
        n8648), .Q(N2985) );
  AO21X1 U8702 ( .IN1(n8419), .IN2(n8633), .IN3(n8422), .Q(n8648) );
  INVX0 U8703 ( .INP(n7677), .ZN(n8422) );
  NAND2X0 U8704 ( .IN1(n7536), .IN2(n7298), .QN(n7677) );
  AO222X1 U8705 ( .IN1(n7686), .IN2(n7684), .IN3(n8635), .IN4(n7599), .IN5(
        n7683), .IN6(n8649), .Q(n8633) );
  NOR3X0 U8706 ( .IN1(n7536), .IN2(n8054), .IN3(n7681), .QN(n8419) );
  INVX0 U8707 ( .INP(n8405), .ZN(n7681) );
  AO222X1 U8708 ( .IN1(n7682), .IN2(n7684), .IN3(n7683), .IN4(n7686), .IN5(
        n8649), .IN6(n7599), .Q(n7691) );
  AO222X1 U8709 ( .IN1(n7688), .IN2(n8650), .IN3(n8434), .IN4(n7687), .IN5(
        n7690), .IN6(n8651), .Q(n7686) );
  AO222X1 U8710 ( .IN1(n8434), .IN2(n7689), .IN3(n7690), .IN4(n7687), .IN5(
        n7688), .IN6(n8651), .Q(n7682) );
  AO222X1 U8711 ( .IN1(n7694), .IN2(n8652), .IN3(n7696), .IN4(n7695), .IN5(
        n7698), .IN6(n8653), .Q(n7687) );
  AO222X1 U8712 ( .IN1(n7696), .IN2(n7699), .IN3(n7698), .IN4(n7695), .IN5(
        n7694), .IN6(n8653), .Q(n7689) );
  AO222X1 U8713 ( .IN1(n7701), .IN2(n8654), .IN3(n7703), .IN4(n7700), .IN5(
        n7705), .IN6(n8655), .Q(n7695) );
  AO222X1 U8714 ( .IN1(n7703), .IN2(n7704), .IN3(n7705), .IN4(n7700), .IN5(
        n7701), .IN6(n8655), .Q(n7699) );
  AO222X1 U8715 ( .IN1(n7709), .IN2(n8656), .IN3(n8501), .IN4(n7708), .IN5(
        n8500), .IN6(n8657), .Q(n7700) );
  AO222X1 U8716 ( .IN1(n8501), .IN2(n7711), .IN3(n8500), .IN4(n7708), .IN5(
        n7709), .IN6(n8657), .Q(n7704) );
  AO222X1 U8717 ( .IN1(n7718), .IN2(n8658), .IN3(n7716), .IN4(n7717), .IN5(
        n7714), .IN6(n8659), .Q(n7708) );
  AO222X1 U8718 ( .IN1(n7716), .IN2(n7713), .IN3(n7714), .IN4(n7717), .IN5(
        n7718), .IN6(n8659), .Q(n7711) );
  AO222X1 U8719 ( .IN1(n7724), .IN2(n8660), .IN3(n7722), .IN4(n7723), .IN5(
        n7720), .IN6(n8661), .Q(n7717) );
  AO222X1 U8720 ( .IN1(n7722), .IN2(n7719), .IN3(n7720), .IN4(n7723), .IN5(
        n7724), .IN6(n8661), .Q(n7713) );
  AO221X1 U8721 ( .IN1(n7726), .IN2(n7732), .IN3(n7730), .IN4(n7727), .IN5(
        n8662), .Q(n7723) );
  AO222X1 U8722 ( .IN1(n7735), .IN2(n7725), .IN3(n8663), .IN4(n7728), .IN5(
        n7733), .IN6(n8664), .Q(n8662) );
  AO221X1 U8723 ( .IN1(n7726), .IN2(n7727), .IN3(n7730), .IN4(n7725), .IN5(
        n8665), .Q(n7719) );
  AO222X1 U8724 ( .IN1(n7735), .IN2(n7731), .IN3(n8663), .IN4(n7733), .IN5(
        n7728), .IN6(n7732), .Q(n8665) );
  AO222X1 U8725 ( .IN1(n7739), .IN2(n7736), .IN3(n7737), .IN4(n7740), .IN5(
        n7741), .IN6(n8666), .Q(n7731) );
  AO222X1 U8726 ( .IN1(n7747), .IN2(n8667), .IN3(n7745), .IN4(n7742), .IN5(
        n7743), .IN6(n7746), .Q(n7736) );
  OAI222X1 U8727 ( .IN1(n7753), .IN2(n8668), .IN3(n7751), .IN4(n7748), .IN5(
        n7749), .IN6(n7752), .QN(n7742) );
  OA222X1 U8728 ( .IN1(n7759), .IN2(n8669), .IN3(n7757), .IN4(n7754), .IN5(
        n7755), .IN6(n7758), .Q(n7748) );
  OA222X1 U8729 ( .IN1(n7764), .IN2(n8670), .IN3(n7664), .IN4(n7760), .IN5(
        n7761), .IN6(n7763), .Q(n7754) );
  OA22X1 U8730 ( .IN1(n7766), .IN2(n4483), .IN3(n7765), .IN4(n4484), .Q(n7760)
         );
  AO222X1 U8731 ( .IN1(n7741), .IN2(n8671), .IN3(n7739), .IN4(n7740), .IN5(
        n7737), .IN6(n8666), .Q(n7725) );
  AO222X1 U8732 ( .IN1(n7747), .IN2(n8672), .IN3(n7745), .IN4(n7746), .IN5(
        n7743), .IN6(n8667), .Q(n7740) );
  AO222X1 U8733 ( .IN1(n7626), .IN2(n8673), .IN3(n7643), .IN4(n8674), .IN5(
        n8647), .IN6(n8675), .Q(n7746) );
  INVX0 U8734 ( .INP(n7752), .ZN(n8674) );
  OA222X1 U8735 ( .IN1(n7759), .IN2(n8676), .IN3(n7757), .IN4(n7758), .IN5(
        n7755), .IN6(n8669), .Q(n7752) );
  OA222X1 U8736 ( .IN1(n7764), .IN2(n8677), .IN3(n7664), .IN4(n7763), .IN5(
        n7761), .IN6(n8670), .Q(n7758) );
  OA22X1 U8737 ( .IN1(n7766), .IN2(n4482), .IN3(n7765), .IN4(n4483), .Q(n7763)
         );
  AND2X1 U8738 ( .IN1(n8566), .IN2(n8254), .Q(n7726) );
  NOR2X0 U8739 ( .IN1(n8405), .IN2(n7536), .QN(n8418) );
  INVX0 U8740 ( .INP(n7874), .ZN(n7536) );
  NAND3X0 U8741 ( .IN1(n3627), .IN2(n7098), .IN3(n3628), .QN(n7874) );
  INVX0 U8742 ( .INP(n7529), .ZN(n7098) );
  NAND3X0 U8743 ( .IN1(n3714), .IN2(n3713), .IN3(n3715), .QN(n7529) );
  AO221X1 U8744 ( .IN1(n8678), .IN2(n8679), .IN3(n8680), .IN4(n7526), .IN5(
        n8681), .Q(n8405) );
  AO21X1 U8745 ( .IN1(n8682), .IN2(n8678), .IN3(n8683), .Q(n8054) );
  AO222X1 U8746 ( .IN1(n8625), .IN2(n7599), .IN3(n7683), .IN4(n8635), .IN5(
        n8649), .IN6(n7684), .Q(n8623) );
  AO222X1 U8747 ( .IN1(n7688), .IN2(n8684), .IN3(n7690), .IN4(n8650), .IN5(
        n8434), .IN6(n8651), .Q(n8649) );
  AO222X1 U8748 ( .IN1(n7696), .IN2(n8653), .IN3(n7698), .IN4(n8652), .IN5(
        n7694), .IN6(n8685), .Q(n8651) );
  AO222X1 U8749 ( .IN1(n7703), .IN2(n8655), .IN3(n7705), .IN4(n8654), .IN5(
        n7701), .IN6(n8686), .Q(n8653) );
  AO222X1 U8750 ( .IN1(n8501), .IN2(n8657), .IN3(n8500), .IN4(n8656), .IN5(
        n7709), .IN6(n8687), .Q(n8655) );
  AO222X1 U8751 ( .IN1(n7716), .IN2(n8659), .IN3(n7714), .IN4(n8658), .IN5(
        n7718), .IN6(n8688), .Q(n8657) );
  AO222X1 U8752 ( .IN1(n7722), .IN2(n8661), .IN3(n7720), .IN4(n8660), .IN5(
        n7724), .IN6(n8689), .Q(n8659) );
  AO221X1 U8753 ( .IN1(n7730), .IN2(n7732), .IN3(n7733), .IN4(n8690), .IN5(
        n8691), .Q(n8661) );
  AO222X1 U8754 ( .IN1(n7735), .IN2(n7727), .IN3(n8663), .IN4(n8566), .IN5(
        n7728), .IN6(n8664), .Q(n8691) );
  AND2X1 U8755 ( .IN1(n8254), .IN2(n8692), .Q(n8663) );
  AO222X1 U8756 ( .IN1(n7741), .IN2(n8693), .IN3(n7739), .IN4(n8666), .IN5(
        n7737), .IN6(n8671), .Q(n7727) );
  AO222X1 U8757 ( .IN1(n7747), .IN2(n8694), .IN3(n7745), .IN4(n8667), .IN5(
        n7743), .IN6(n8672), .Q(n8666) );
  AO222X1 U8758 ( .IN1(n7626), .IN2(n8695), .IN3(n7643), .IN4(n8675), .IN5(
        n8647), .IN6(n8673), .Q(n8667) );
  INVX0 U8759 ( .INP(n8668), .ZN(n8675) );
  OA222X1 U8760 ( .IN1(n7759), .IN2(n8696), .IN3(n7757), .IN4(n8669), .IN5(
        n7755), .IN6(n8676), .Q(n8668) );
  INVX0 U8761 ( .INP(n8697), .ZN(n7755) );
  OA222X1 U8762 ( .IN1(n7764), .IN2(n8698), .IN3(n7664), .IN4(n8670), .IN5(
        n7761), .IN6(n8677), .Q(n8669) );
  OA22X1 U8763 ( .IN1(n7766), .IN2(n4481), .IN3(n7765), .IN4(n4482), .Q(n8670)
         );
  INVX0 U8764 ( .INP(n8699), .ZN(n7759) );
  AO222X1 U8765 ( .IN1(n8434), .IN2(n8650), .IN3(n7688), .IN4(n8636), .IN5(
        n7690), .IN6(n8684), .Q(n8635) );
  AO222X1 U8766 ( .IN1(n7696), .IN2(n8652), .IN3(n7694), .IN4(n8700), .IN5(
        n7698), .IN6(n8685), .Q(n8650) );
  AO222X1 U8767 ( .IN1(n7701), .IN2(n8701), .IN3(n7703), .IN4(n8654), .IN5(
        n7705), .IN6(n8686), .Q(n8652) );
  AO222X1 U8768 ( .IN1(n7709), .IN2(n8702), .IN3(n8501), .IN4(n8656), .IN5(
        n8500), .IN6(n8687), .Q(n8654) );
  AO222X1 U8769 ( .IN1(n7718), .IN2(n8703), .IN3(n7716), .IN4(n8658), .IN5(
        n7714), .IN6(n8688), .Q(n8656) );
  AO222X1 U8770 ( .IN1(n7724), .IN2(n8704), .IN3(n7722), .IN4(n8660), .IN5(
        n7720), .IN6(n8689), .Q(n8658) );
  AO221X1 U8771 ( .IN1(n7733), .IN2(n8705), .IN3(n7728), .IN4(n8690), .IN5(
        n8706), .Q(n8660) );
  AO22X1 U8772 ( .IN1(n8566), .IN2(n8664), .IN3(n7735), .IN4(n7732), .Q(n8706)
         );
  AO222X1 U8773 ( .IN1(n7741), .IN2(n8707), .IN3(n7739), .IN4(n8671), .IN5(
        n7737), .IN6(n8693), .Q(n7732) );
  AO222X1 U8774 ( .IN1(n7747), .IN2(n8708), .IN3(n7745), .IN4(n8672), .IN5(
        n7743), .IN6(n8694), .Q(n8671) );
  AO222X1 U8775 ( .IN1(n7626), .IN2(n8709), .IN3(n7643), .IN4(n8673), .IN5(
        n8647), .IN6(n8695), .Q(n8672) );
  AO222X1 U8776 ( .IN1(n8699), .IN2(n8710), .IN3(n8711), .IN4(n8712), .IN5(
        n8697), .IN6(n8713), .Q(n8673) );
  INVX0 U8777 ( .INP(n8676), .ZN(n8712) );
  OA222X1 U8778 ( .IN1(n7764), .IN2(n8714), .IN3(n7664), .IN4(n8677), .IN5(
        n7761), .IN6(n8698), .Q(n8676) );
  OA22X1 U8779 ( .IN1(n7766), .IN2(n4480), .IN3(n7765), .IN4(n4481), .Q(n8677)
         );
  AND2X1 U8780 ( .IN1(n8566), .IN2(n8099), .Q(n7735) );
  AO22X1 U8781 ( .IN1(n7730), .IN2(n8692), .IN3(n8254), .IN4(n8715), .Q(n8664)
         );
  NOR2X0 U8782 ( .IN1(n7684), .IN2(n7599), .QN(n7683) );
  INVX0 U8783 ( .INP(n7606), .ZN(n7684) );
  NAND2X0 U8784 ( .IN1(n8716), .IN2(n8717), .QN(n7606) );
  AO21X1 U8785 ( .IN1(n8682), .IN2(n8718), .IN3(n8719), .Q(n7599) );
  AO222X1 U8786 ( .IN1(n7688), .IN2(n8626), .IN3(n7690), .IN4(n8636), .IN5(
        n8434), .IN6(n8684), .Q(n8625) );
  AO222X1 U8787 ( .IN1(n7694), .IN2(n8720), .IN3(n7698), .IN4(n8700), .IN5(
        n7696), .IN6(n8685), .Q(n8684) );
  AO222X1 U8788 ( .IN1(n7701), .IN2(n8721), .IN3(n7705), .IN4(n8701), .IN5(
        n7703), .IN6(n8686), .Q(n8685) );
  AO222X1 U8789 ( .IN1(n7709), .IN2(n8722), .IN3(n8500), .IN4(n8702), .IN5(
        n8501), .IN6(n8687), .Q(n8686) );
  AO222X1 U8790 ( .IN1(n7718), .IN2(n8723), .IN3(n7714), .IN4(n8703), .IN5(
        n7716), .IN6(n8688), .Q(n8687) );
  AO222X1 U8791 ( .IN1(n7724), .IN2(n8724), .IN3(n7720), .IN4(n8704), .IN5(
        n7722), .IN6(n8689), .Q(n8688) );
  AO222X1 U8792 ( .IN1(n8566), .IN2(n8690), .IN3(n7728), .IN4(n8705), .IN5(
        n7733), .IN6(n8725), .Q(n8689) );
  AO222X1 U8793 ( .IN1(n8099), .IN2(n8692), .IN3(n7730), .IN4(n8715), .IN5(
        n8726), .IN6(n8254), .Q(n8690) );
  AO222X1 U8794 ( .IN1(n7741), .IN2(n8727), .IN3(n7739), .IN4(n8693), .IN5(
        n7737), .IN6(n8707), .Q(n8692) );
  AO222X1 U8795 ( .IN1(n7747), .IN2(n8728), .IN3(n7745), .IN4(n8694), .IN5(
        n7743), .IN6(n8708), .Q(n8693) );
  AO222X1 U8796 ( .IN1(n7626), .IN2(n8729), .IN3(n7643), .IN4(n8695), .IN5(
        n8647), .IN6(n8709), .Q(n8694) );
  AO222X1 U8797 ( .IN1(n8699), .IN2(n8730), .IN3(n8711), .IN4(n8713), .IN5(
        n8697), .IN6(n8710), .Q(n8695) );
  INVX0 U8798 ( .INP(n8696), .ZN(n8713) );
  OA222X1 U8799 ( .IN1(n7764), .IN2(n8731), .IN3(n7664), .IN4(n8698), .IN5(
        n7761), .IN6(n8714), .Q(n8696) );
  OA22X1 U8800 ( .IN1(n7766), .IN2(n4479), .IN3(n7765), .IN4(n4480), .Q(n8698)
         );
  INVX0 U8801 ( .INP(n8525), .ZN(n7664) );
  NOR2X0 U8802 ( .IN1(n8406), .IN2(n8338), .QN(n8434) );
  AO222X1 U8803 ( .IN1(n7696), .IN2(n8700), .IN3(n7694), .IN4(n8637), .IN5(
        n7698), .IN6(n8720), .Q(n8636) );
  AO222X1 U8804 ( .IN1(n7703), .IN2(n8701), .IN3(n7701), .IN4(n8732), .IN5(
        n7705), .IN6(n8721), .Q(n8700) );
  AO222X1 U8805 ( .IN1(n8501), .IN2(n8702), .IN3(n7709), .IN4(n8733), .IN5(
        n8500), .IN6(n8722), .Q(n8701) );
  AO222X1 U8806 ( .IN1(n7716), .IN2(n8703), .IN3(n7718), .IN4(n8734), .IN5(
        n7714), .IN6(n8723), .Q(n8702) );
  AO222X1 U8807 ( .IN1(n7722), .IN2(n8704), .IN3(n7724), .IN4(n8735), .IN5(
        n7720), .IN6(n8724), .Q(n8703) );
  AO222X1 U8808 ( .IN1(n8566), .IN2(n8705), .IN3(n7733), .IN4(n8736), .IN5(
        n7728), .IN6(n8725), .Q(n8704) );
  AO222X1 U8809 ( .IN1(n8737), .IN2(n8254), .IN3(n8099), .IN4(n8715), .IN5(
        n7730), .IN6(n8726), .Q(n8705) );
  AO222X1 U8810 ( .IN1(n7737), .IN2(n8727), .IN3(n7739), .IN4(n8707), .IN5(
        n7741), .IN6(n8738), .Q(n8715) );
  AO222X1 U8811 ( .IN1(n7743), .IN2(n8728), .IN3(n7745), .IN4(n8708), .IN5(
        n7747), .IN6(n8739), .Q(n8707) );
  AO222X1 U8812 ( .IN1(n8647), .IN2(n8729), .IN3(n7643), .IN4(n8709), .IN5(
        n7626), .IN6(n8740), .Q(n8708) );
  AO222X1 U8813 ( .IN1(n8697), .IN2(n8730), .IN3(n8711), .IN4(n8710), .IN5(
        n8699), .IN6(n8741), .Q(n8709) );
  AO222X1 U8814 ( .IN1(n8536), .IN2(n8742), .IN3(n8525), .IN4(n8743), .IN5(
        n8538), .IN6(n8744), .Q(n8710) );
  INVX0 U8815 ( .INP(n8714), .ZN(n8743) );
  OA22X1 U8816 ( .IN1(n7766), .IN2(n4478), .IN3(n7765), .IN4(n4479), .Q(n8714)
         );
  XOR2X1 U8817 ( .IN1(n8406), .IN2(n8338), .Q(n7690) );
  AO222X1 U8818 ( .IN1(n7694), .IN2(n8627), .IN3(n7698), .IN4(n8637), .IN5(
        n7696), .IN6(n8720), .Q(n8626) );
  AO222X1 U8819 ( .IN1(n7701), .IN2(n8745), .IN3(n7705), .IN4(n8732), .IN5(
        n7703), .IN6(n8721), .Q(n8720) );
  AO222X1 U8820 ( .IN1(n7709), .IN2(n8746), .IN3(n8500), .IN4(n8733), .IN5(
        n8501), .IN6(n8722), .Q(n8721) );
  AO222X1 U8821 ( .IN1(n7718), .IN2(n8747), .IN3(n7714), .IN4(n8734), .IN5(
        n7716), .IN6(n8723), .Q(n8722) );
  AO222X1 U8822 ( .IN1(n7724), .IN2(n8748), .IN3(n7720), .IN4(n8735), .IN5(
        n7722), .IN6(n8724), .Q(n8723) );
  AO222X1 U8823 ( .IN1(n7733), .IN2(n8749), .IN3(n7728), .IN4(n8736), .IN5(
        n8566), .IN6(n8725), .Q(n8724) );
  AO222X1 U8824 ( .IN1(n8750), .IN2(n8254), .IN3(n7730), .IN4(n8737), .IN5(
        n8099), .IN6(n8726), .Q(n8725) );
  AO222X1 U8825 ( .IN1(n7741), .IN2(n8751), .IN3(n7737), .IN4(n8738), .IN5(
        n7739), .IN6(n8727), .Q(n8726) );
  AO222X1 U8826 ( .IN1(n7747), .IN2(n8752), .IN3(n7745), .IN4(n8728), .IN5(
        n7743), .IN6(n8739), .Q(n8727) );
  AO222X1 U8827 ( .IN1(n8753), .IN2(n7626), .IN3(n7643), .IN4(n8729), .IN5(
        n8647), .IN6(n8740), .Q(n8728) );
  AO222X1 U8828 ( .IN1(n8699), .IN2(n8754), .IN3(n8711), .IN4(n8730), .IN5(
        n8697), .IN6(n8741), .Q(n8729) );
  AO222X1 U8829 ( .IN1(n8538), .IN2(n8755), .IN3(n8525), .IN4(n8742), .IN5(
        n8536), .IN6(n8744), .Q(n8730) );
  INVX0 U8830 ( .INP(n8731), .ZN(n8742) );
  OA22X1 U8831 ( .IN1(n7766), .IN2(n4477), .IN3(n7765), .IN4(n4478), .Q(n8731)
         );
  NOR2X0 U8832 ( .IN1(n8337), .IN2(n8253), .QN(n7696) );
  AO222X1 U8833 ( .IN1(n7703), .IN2(n8732), .IN3(n7701), .IN4(n8638), .IN5(
        n7705), .IN6(n8745), .Q(n8637) );
  AO222X1 U8834 ( .IN1(n8501), .IN2(n8733), .IN3(n7709), .IN4(n8756), .IN5(
        n8500), .IN6(n8746), .Q(n8732) );
  AO222X1 U8835 ( .IN1(n7716), .IN2(n8734), .IN3(n7718), .IN4(n8757), .IN5(
        n7714), .IN6(n8747), .Q(n8733) );
  AO222X1 U8836 ( .IN1(n7722), .IN2(n8735), .IN3(n7724), .IN4(n8758), .IN5(
        n7720), .IN6(n8748), .Q(n8734) );
  AO222X1 U8837 ( .IN1(n8566), .IN2(n8736), .IN3(n7733), .IN4(n8759), .IN5(
        n7728), .IN6(n8749), .Q(n8735) );
  AO222X1 U8838 ( .IN1(n8099), .IN2(n8737), .IN3(n8760), .IN4(n8254), .IN5(
        n7730), .IN6(n8750), .Q(n8736) );
  AO222X1 U8839 ( .IN1(n7739), .IN2(n8738), .IN3(n7741), .IN4(n8761), .IN5(
        n7737), .IN6(n8751), .Q(n8737) );
  AO222X1 U8840 ( .IN1(n7747), .IN2(n8762), .IN3(n7745), .IN4(n8739), .IN5(
        n7743), .IN6(n8752), .Q(n8738) );
  AO222X1 U8841 ( .IN1(n8763), .IN2(n7626), .IN3(n7643), .IN4(n8740), .IN5(
        n8647), .IN6(n8753), .Q(n8739) );
  AO222X1 U8842 ( .IN1(n8699), .IN2(n8764), .IN3(n8711), .IN4(n8741), .IN5(
        n8697), .IN6(n8754), .Q(n8740) );
  AO222X1 U8843 ( .IN1(n8538), .IN2(n8765), .IN3(n8525), .IN4(n8744), .IN5(
        n8536), .IN6(n8755), .Q(n8741) );
  AO22X1 U8844 ( .IN1(n8766), .IN2(n7276), .IN3(n8767), .IN4(n7275), .Q(n8744)
         );
  XOR2X1 U8845 ( .IN1(n8337), .IN2(n8253), .Q(n7698) );
  INVX0 U8846 ( .INP(n8768), .ZN(n8253) );
  AO222X1 U8847 ( .IN1(n7701), .IN2(n8628), .IN3(n7705), .IN4(n8638), .IN5(
        n7703), .IN6(n8745), .Q(n8627) );
  AO222X1 U8848 ( .IN1(n7709), .IN2(n8769), .IN3(n8500), .IN4(n8756), .IN5(
        n8501), .IN6(n8746), .Q(n8745) );
  AO222X1 U8849 ( .IN1(n7718), .IN2(n8770), .IN3(n7714), .IN4(n8757), .IN5(
        n7716), .IN6(n8747), .Q(n8746) );
  AO222X1 U8850 ( .IN1(n7724), .IN2(n8771), .IN3(n7720), .IN4(n8758), .IN5(
        n7722), .IN6(n8748), .Q(n8747) );
  AO222X1 U8851 ( .IN1(n7733), .IN2(n8772), .IN3(n7728), .IN4(n8759), .IN5(
        n8566), .IN6(n8749), .Q(n8748) );
  AO222X1 U8852 ( .IN1(n8773), .IN2(n8254), .IN3(n7730), .IN4(n8760), .IN5(
        n8099), .IN6(n8750), .Q(n8749) );
  AO222X1 U8853 ( .IN1(n7741), .IN2(n8774), .IN3(n7737), .IN4(n8761), .IN5(
        n7739), .IN6(n8751), .Q(n8750) );
  AO222X1 U8854 ( .IN1(n7747), .IN2(n8775), .IN3(n7743), .IN4(n8762), .IN5(
        n7745), .IN6(n8752), .Q(n8751) );
  AO222X1 U8855 ( .IN1(n8776), .IN2(n7626), .IN3(n8647), .IN4(n8763), .IN5(
        n7643), .IN6(n8753), .Q(n8752) );
  AO222X1 U8856 ( .IN1(n8699), .IN2(n8777), .IN3(n8697), .IN4(n8764), .IN5(
        n8711), .IN6(n8754), .Q(n8753) );
  AO222X1 U8857 ( .IN1(n8538), .IN2(n8778), .IN3(n8536), .IN4(n8765), .IN5(
        n8525), .IN6(n8755), .Q(n8754) );
  AO222X1 U8858 ( .IN1(n8767), .IN2(n7276), .IN3(n8779), .IN4(n7275), .IN5(
        n8766), .IN6(n7277), .Q(n8755) );
  INVX0 U8859 ( .INP(n4477), .ZN(n7275) );
  NOR2X0 U8860 ( .IN1(n8227), .IN2(n7638), .QN(n7703) );
  AO222X1 U8861 ( .IN1(n8501), .IN2(n8756), .IN3(n7709), .IN4(n8639), .IN5(
        n8500), .IN6(n8769), .Q(n8638) );
  AO222X1 U8862 ( .IN1(n7716), .IN2(n8757), .IN3(n7718), .IN4(n8780), .IN5(
        n7714), .IN6(n8770), .Q(n8756) );
  AO222X1 U8863 ( .IN1(n7722), .IN2(n8758), .IN3(n7724), .IN4(n8781), .IN5(
        n7720), .IN6(n8771), .Q(n8757) );
  AO222X1 U8864 ( .IN1(n8566), .IN2(n8759), .IN3(n7733), .IN4(n8782), .IN5(
        n7728), .IN6(n8772), .Q(n8758) );
  AO222X1 U8865 ( .IN1(n8099), .IN2(n8760), .IN3(n8783), .IN4(n8254), .IN5(
        n7730), .IN6(n8773), .Q(n8759) );
  AO222X1 U8866 ( .IN1(n7739), .IN2(n8761), .IN3(n7741), .IN4(n8784), .IN5(
        n7737), .IN6(n8774), .Q(n8760) );
  AO222X1 U8867 ( .IN1(n7745), .IN2(n8762), .IN3(n7747), .IN4(n8785), .IN5(
        n7743), .IN6(n8775), .Q(n8761) );
  AO222X1 U8868 ( .IN1(n7643), .IN2(n8763), .IN3(n8786), .IN4(n7626), .IN5(
        n8647), .IN6(n8776), .Q(n8762) );
  AO222X1 U8869 ( .IN1(n8711), .IN2(n8764), .IN3(n8699), .IN4(n8787), .IN5(
        n8697), .IN6(n8777), .Q(n8763) );
  AO222X1 U8870 ( .IN1(n8525), .IN2(n8765), .IN3(n8538), .IN4(n8788), .IN5(
        n8536), .IN6(n8778), .Q(n8764) );
  AO222X1 U8871 ( .IN1(n8767), .IN2(n7277), .IN3(n8779), .IN4(n7276), .IN5(
        n8766), .IN6(n7278), .Q(n8765) );
  INVX0 U8872 ( .INP(n4476), .ZN(n7276) );
  XOR2X1 U8873 ( .IN1(n8227), .IN2(n7638), .Q(n7705) );
  AO222X1 U8874 ( .IN1(n7709), .IN2(n8629), .IN3(n8500), .IN4(n8639), .IN5(
        n8501), .IN6(n8769), .Q(n8628) );
  AO222X1 U8875 ( .IN1(n7718), .IN2(n8789), .IN3(n7714), .IN4(n8780), .IN5(
        n7716), .IN6(n8770), .Q(n8769) );
  AO222X1 U8876 ( .IN1(n7724), .IN2(n8790), .IN3(n7720), .IN4(n8781), .IN5(
        n7722), .IN6(n8771), .Q(n8770) );
  AO222X1 U8877 ( .IN1(n7733), .IN2(n8791), .IN3(n7728), .IN4(n8782), .IN5(
        n8566), .IN6(n8772), .Q(n8771) );
  AO222X1 U8878 ( .IN1(n8792), .IN2(n8254), .IN3(n7730), .IN4(n8783), .IN5(
        n8099), .IN6(n8773), .Q(n8772) );
  AO222X1 U8879 ( .IN1(n7741), .IN2(n8793), .IN3(n7737), .IN4(n8784), .IN5(
        n7739), .IN6(n8774), .Q(n8773) );
  AO222X1 U8880 ( .IN1(n7747), .IN2(n8794), .IN3(n7743), .IN4(n8785), .IN5(
        n7745), .IN6(n8775), .Q(n8774) );
  AO222X1 U8881 ( .IN1(n8795), .IN2(n7626), .IN3(n8647), .IN4(n8786), .IN5(
        n7643), .IN6(n8776), .Q(n8775) );
  AO222X1 U8882 ( .IN1(n8699), .IN2(n8796), .IN3(n8697), .IN4(n8787), .IN5(
        n8711), .IN6(n8777), .Q(n8776) );
  AO222X1 U8883 ( .IN1(n8538), .IN2(n8797), .IN3(n8536), .IN4(n8788), .IN5(
        n8525), .IN6(n8778), .Q(n8777) );
  AO222X1 U8884 ( .IN1(n8767), .IN2(n7278), .IN3(n8779), .IN4(n7277), .IN5(
        n8766), .IN6(n7279), .Q(n8778) );
  INVX0 U8885 ( .INP(n4475), .ZN(n7277) );
  NOR2X0 U8886 ( .IN1(n8319), .IN2(n7712), .QN(n8501) );
  INVX0 U8887 ( .INP(n7706), .ZN(n8319) );
  AO222X1 U8888 ( .IN1(n7716), .IN2(n8780), .IN3(n7718), .IN4(n8640), .IN5(
        n7714), .IN6(n8789), .Q(n8639) );
  AO222X1 U8889 ( .IN1(n7722), .IN2(n8781), .IN3(n7724), .IN4(n8798), .IN5(
        n7720), .IN6(n8790), .Q(n8780) );
  AO222X1 U8890 ( .IN1(n8566), .IN2(n8782), .IN3(n7733), .IN4(n8799), .IN5(
        n7728), .IN6(n8791), .Q(n8781) );
  AO222X1 U8891 ( .IN1(n8099), .IN2(n8783), .IN3(n8800), .IN4(n8254), .IN5(
        n7730), .IN6(n8792), .Q(n8782) );
  AO222X1 U8892 ( .IN1(n7739), .IN2(n8784), .IN3(n7741), .IN4(n8801), .IN5(
        n7737), .IN6(n8793), .Q(n8783) );
  AO222X1 U8893 ( .IN1(n7745), .IN2(n8785), .IN3(n7747), .IN4(n8802), .IN5(
        n7743), .IN6(n8794), .Q(n8784) );
  AO222X1 U8894 ( .IN1(n7643), .IN2(n8786), .IN3(n8803), .IN4(n7626), .IN5(
        n8647), .IN6(n8795), .Q(n8785) );
  AO222X1 U8895 ( .IN1(n8711), .IN2(n8787), .IN3(n8699), .IN4(n8804), .IN5(
        n8697), .IN6(n8796), .Q(n8786) );
  AO222X1 U8896 ( .IN1(n8525), .IN2(n8788), .IN3(n8538), .IN4(n8805), .IN5(
        n8536), .IN6(n8797), .Q(n8787) );
  AO222X1 U8897 ( .IN1(n8767), .IN2(n7279), .IN3(n8779), .IN4(n7278), .IN5(
        n8766), .IN6(n7280), .Q(n8788) );
  INVX0 U8898 ( .INP(n4474), .ZN(n7278) );
  XOR2X1 U8899 ( .IN1(n8806), .IN2(n7706), .Q(n8500) );
  AO222X1 U8900 ( .IN1(n7718), .IN2(n8630), .IN3(n7714), .IN4(n8640), .IN5(
        n7716), .IN6(n8789), .Q(n8629) );
  AO222X1 U8901 ( .IN1(n7724), .IN2(n8807), .IN3(n7720), .IN4(n8798), .IN5(
        n7722), .IN6(n8790), .Q(n8789) );
  AO222X1 U8902 ( .IN1(n7733), .IN2(n8808), .IN3(n7728), .IN4(n8799), .IN5(
        n8566), .IN6(n8791), .Q(n8790) );
  AO222X1 U8903 ( .IN1(n8809), .IN2(n8254), .IN3(n7730), .IN4(n8800), .IN5(
        n8099), .IN6(n8792), .Q(n8791) );
  AO222X1 U8904 ( .IN1(n7741), .IN2(n8810), .IN3(n7737), .IN4(n8801), .IN5(
        n7739), .IN6(n8793), .Q(n8792) );
  AO222X1 U8905 ( .IN1(n7747), .IN2(n8811), .IN3(n7743), .IN4(n8802), .IN5(
        n7745), .IN6(n8794), .Q(n8793) );
  AO222X1 U8906 ( .IN1(n8812), .IN2(n7626), .IN3(n8647), .IN4(n8803), .IN5(
        n7643), .IN6(n8795), .Q(n8794) );
  AO222X1 U8907 ( .IN1(n8699), .IN2(n8813), .IN3(n8697), .IN4(n8804), .IN5(
        n8711), .IN6(n8796), .Q(n8795) );
  AO222X1 U8908 ( .IN1(n8538), .IN2(n8814), .IN3(n8536), .IN4(n8805), .IN5(
        n8525), .IN6(n8797), .Q(n8796) );
  AO222X1 U8909 ( .IN1(n8767), .IN2(n7280), .IN3(n8779), .IN4(n7279), .IN5(
        n8766), .IN6(n7281), .Q(n8797) );
  INVX0 U8910 ( .INP(n4473), .ZN(n7279) );
  NOR2X0 U8911 ( .IN1(n8391), .IN2(n7671), .QN(n7716) );
  AO222X1 U8912 ( .IN1(n7722), .IN2(n8798), .IN3(n7724), .IN4(n8641), .IN5(
        n7720), .IN6(n8807), .Q(n8640) );
  AO222X1 U8913 ( .IN1(n8566), .IN2(n8799), .IN3(n7733), .IN4(n8815), .IN5(
        n7728), .IN6(n8808), .Q(n8798) );
  AO222X1 U8914 ( .IN1(n8099), .IN2(n8800), .IN3(n8816), .IN4(n8254), .IN5(
        n7730), .IN6(n8809), .Q(n8799) );
  AO222X1 U8915 ( .IN1(n7739), .IN2(n8801), .IN3(n7741), .IN4(n8817), .IN5(
        n7737), .IN6(n8810), .Q(n8800) );
  AO222X1 U8916 ( .IN1(n7745), .IN2(n8802), .IN3(n7747), .IN4(n8818), .IN5(
        n7743), .IN6(n8811), .Q(n8801) );
  AO222X1 U8917 ( .IN1(n7643), .IN2(n8803), .IN3(n8819), .IN4(n7626), .IN5(
        n8647), .IN6(n8812), .Q(n8802) );
  AO222X1 U8918 ( .IN1(n8711), .IN2(n8804), .IN3(n8699), .IN4(n8820), .IN5(
        n8697), .IN6(n8813), .Q(n8803) );
  AO222X1 U8919 ( .IN1(n8525), .IN2(n8805), .IN3(n8538), .IN4(n8821), .IN5(
        n8536), .IN6(n8814), .Q(n8804) );
  AO222X1 U8920 ( .IN1(n8767), .IN2(n7281), .IN3(n8779), .IN4(n7280), .IN5(
        n8766), .IN6(n7282), .Q(n8805) );
  INVX0 U8921 ( .INP(n4472), .ZN(n7280) );
  XOR2X1 U8922 ( .IN1(n7671), .IN2(n8391), .Q(n7714) );
  AO222X1 U8923 ( .IN1(n7724), .IN2(n8631), .IN3(n7720), .IN4(n8641), .IN5(
        n7722), .IN6(n8807), .Q(n8630) );
  AO222X1 U8924 ( .IN1(n7733), .IN2(n8822), .IN3(n7728), .IN4(n8815), .IN5(
        n8566), .IN6(n8808), .Q(n8807) );
  AO222X1 U8925 ( .IN1(n8823), .IN2(n8254), .IN3(n7730), .IN4(n8816), .IN5(
        n8099), .IN6(n8809), .Q(n8808) );
  AO222X1 U8926 ( .IN1(n7741), .IN2(n8824), .IN3(n7737), .IN4(n8817), .IN5(
        n7739), .IN6(n8810), .Q(n8809) );
  AO222X1 U8927 ( .IN1(n7747), .IN2(n8825), .IN3(n7743), .IN4(n8818), .IN5(
        n7745), .IN6(n8811), .Q(n8810) );
  AO222X1 U8928 ( .IN1(n8826), .IN2(n7626), .IN3(n8647), .IN4(n8819), .IN5(
        n7643), .IN6(n8812), .Q(n8811) );
  AO222X1 U8929 ( .IN1(n8699), .IN2(n8827), .IN3(n8697), .IN4(n8820), .IN5(
        n8711), .IN6(n8813), .Q(n8812) );
  AO222X1 U8930 ( .IN1(n8538), .IN2(n8828), .IN3(n8536), .IN4(n8821), .IN5(
        n8525), .IN6(n8814), .Q(n8813) );
  AO222X1 U8931 ( .IN1(n8767), .IN2(n7282), .IN3(n8779), .IN4(n7281), .IN5(
        n8766), .IN6(n7283), .Q(n8814) );
  INVX0 U8932 ( .INP(n4471), .ZN(n7281) );
  NOR2X0 U8933 ( .IN1(n8318), .IN2(n7644), .QN(n7722) );
  AO222X1 U8934 ( .IN1(n8566), .IN2(n8815), .IN3(n7733), .IN4(n8642), .IN5(
        n7728), .IN6(n8822), .Q(n8641) );
  AO222X1 U8935 ( .IN1(n8099), .IN2(n8816), .IN3(n8829), .IN4(n8254), .IN5(
        n7730), .IN6(n8823), .Q(n8815) );
  AO222X1 U8936 ( .IN1(n7739), .IN2(n8817), .IN3(n7741), .IN4(n8830), .IN5(
        n7737), .IN6(n8824), .Q(n8816) );
  AO222X1 U8937 ( .IN1(n7745), .IN2(n8818), .IN3(n7747), .IN4(n8831), .IN5(
        n7743), .IN6(n8825), .Q(n8817) );
  AO222X1 U8938 ( .IN1(n7643), .IN2(n8819), .IN3(n8832), .IN4(n7626), .IN5(
        n8647), .IN6(n8826), .Q(n8818) );
  AO222X1 U8939 ( .IN1(n8711), .IN2(n8820), .IN3(n8699), .IN4(n8833), .IN5(
        n8697), .IN6(n8827), .Q(n8819) );
  AO222X1 U8940 ( .IN1(n8525), .IN2(n8821), .IN3(n8538), .IN4(n8834), .IN5(
        n8536), .IN6(n8828), .Q(n8820) );
  AO222X1 U8941 ( .IN1(n8767), .IN2(n7283), .IN3(n8779), .IN4(n7282), .IN5(
        n8766), .IN6(n7284), .Q(n8821) );
  INVX0 U8942 ( .INP(n4470), .ZN(n7282) );
  XOR2X1 U8943 ( .IN1(n8318), .IN2(n7644), .Q(n7720) );
  AO222X1 U8944 ( .IN1(n7733), .IN2(n8632), .IN3(n7728), .IN4(n8642), .IN5(
        n8566), .IN6(n8822), .Q(n8631) );
  AO222X1 U8945 ( .IN1(n8835), .IN2(n8254), .IN3(n7730), .IN4(n8829), .IN5(
        n8099), .IN6(n8823), .Q(n8822) );
  AO222X1 U8946 ( .IN1(n7741), .IN2(n8836), .IN3(n7737), .IN4(n8830), .IN5(
        n7739), .IN6(n8824), .Q(n8823) );
  AO222X1 U8947 ( .IN1(n7747), .IN2(n8837), .IN3(n7743), .IN4(n8831), .IN5(
        n7745), .IN6(n8825), .Q(n8824) );
  AO222X1 U8948 ( .IN1(n8838), .IN2(n7626), .IN3(n8647), .IN4(n8832), .IN5(
        n7643), .IN6(n8826), .Q(n8825) );
  AO222X1 U8949 ( .IN1(n8699), .IN2(n8839), .IN3(n8697), .IN4(n8833), .IN5(
        n8711), .IN6(n8827), .Q(n8826) );
  AO222X1 U8950 ( .IN1(n8538), .IN2(n8840), .IN3(n8536), .IN4(n8834), .IN5(
        n8525), .IN6(n8828), .Q(n8827) );
  AO222X1 U8951 ( .IN1(n8767), .IN2(n7284), .IN3(n8779), .IN4(n7283), .IN5(
        n8766), .IN6(n7285), .Q(n8828) );
  INVX0 U8952 ( .INP(n4469), .ZN(n7283) );
  NOR2X0 U8953 ( .IN1(n8053), .IN2(n7650), .QN(n8566) );
  AO222X1 U8954 ( .IN1(n8099), .IN2(n8829), .IN3(n8643), .IN4(n8254), .IN5(
        n7730), .IN6(n8835), .Q(n8642) );
  AO222X1 U8955 ( .IN1(n7739), .IN2(n8830), .IN3(n7741), .IN4(n8841), .IN5(
        n7737), .IN6(n8836), .Q(n8829) );
  AO222X1 U8956 ( .IN1(n7745), .IN2(n8831), .IN3(n7747), .IN4(n8842), .IN5(
        n7743), .IN6(n8837), .Q(n8830) );
  AO222X1 U8957 ( .IN1(n7643), .IN2(n8832), .IN3(n8843), .IN4(n7626), .IN5(
        n8647), .IN6(n8838), .Q(n8831) );
  AO222X1 U8958 ( .IN1(n8711), .IN2(n8833), .IN3(n8699), .IN4(n8844), .IN5(
        n8697), .IN6(n8839), .Q(n8832) );
  AO222X1 U8959 ( .IN1(n8525), .IN2(n8834), .IN3(n8538), .IN4(n8845), .IN5(
        n8536), .IN6(n8840), .Q(n8833) );
  AO222X1 U8960 ( .IN1(n8767), .IN2(n7285), .IN3(n8779), .IN4(n7284), .IN5(
        n8766), .IN6(n7286), .Q(n8834) );
  INVX0 U8961 ( .INP(n4468), .ZN(n7284) );
  XOR2X1 U8962 ( .IN1(n8053), .IN2(n7650), .Q(n7728) );
  AO222X1 U8963 ( .IN1(n8610), .IN2(n8254), .IN3(n7730), .IN4(n8643), .IN5(
        n8099), .IN6(n8835), .Q(n8632) );
  AO222X1 U8964 ( .IN1(n7741), .IN2(n8846), .IN3(n7737), .IN4(n8841), .IN5(
        n7739), .IN6(n8836), .Q(n8835) );
  AO222X1 U8965 ( .IN1(n7747), .IN2(n8847), .IN3(n7743), .IN4(n8842), .IN5(
        n7745), .IN6(n8837), .Q(n8836) );
  AO222X1 U8966 ( .IN1(n8848), .IN2(n7626), .IN3(n8647), .IN4(n8843), .IN5(
        n7643), .IN6(n8838), .Q(n8837) );
  AO222X1 U8967 ( .IN1(n8699), .IN2(n8849), .IN3(n8697), .IN4(n8844), .IN5(
        n8711), .IN6(n8839), .Q(n8838) );
  AO222X1 U8968 ( .IN1(n8538), .IN2(n8850), .IN3(n8536), .IN4(n8845), .IN5(
        n8525), .IN6(n8840), .Q(n8839) );
  AO222X1 U8969 ( .IN1(n8767), .IN2(n7286), .IN3(n8779), .IN4(n7285), .IN5(
        n8766), .IN6(n7287), .Q(n8840) );
  INVX0 U8970 ( .INP(n4467), .ZN(n7285) );
  AO222X1 U8971 ( .IN1(n7739), .IN2(n8841), .IN3(n7741), .IN4(n8644), .IN5(
        n7737), .IN6(n8846), .Q(n8643) );
  AO222X1 U8972 ( .IN1(n7745), .IN2(n8842), .IN3(n7747), .IN4(n8851), .IN5(
        n7743), .IN6(n8847), .Q(n8841) );
  AO222X1 U8973 ( .IN1(n7643), .IN2(n8843), .IN3(n8852), .IN4(n7626), .IN5(
        n8647), .IN6(n8848), .Q(n8842) );
  AO222X1 U8974 ( .IN1(n8711), .IN2(n8844), .IN3(n8699), .IN4(n8853), .IN5(
        n8697), .IN6(n8849), .Q(n8843) );
  AO222X1 U8975 ( .IN1(n8525), .IN2(n8845), .IN3(n8538), .IN4(n8854), .IN5(
        n8536), .IN6(n8850), .Q(n8844) );
  AO222X1 U8976 ( .IN1(n8767), .IN2(n7287), .IN3(n8779), .IN4(n7286), .IN5(
        n8766), .IN6(n7288), .Q(n8845) );
  INVX0 U8977 ( .INP(n4466), .ZN(n7286) );
  NOR2X0 U8978 ( .IN1(n8254), .IN2(n8099), .QN(n7730) );
  INVX0 U8979 ( .INP(n7603), .ZN(n8099) );
  AO221X1 U8980 ( .IN1(n8855), .IN2(n8856), .IN3(n8857), .IN4(n8680), .IN5(
        n8858), .Q(n7603) );
  AO221X1 U8981 ( .IN1(n8855), .IN2(n8859), .IN3(n8679), .IN4(n8860), .IN5(
        n8858), .Q(n8254) );
  INVX0 U8982 ( .INP(n8861), .ZN(n8858) );
  AO222X1 U8983 ( .IN1(n7741), .IN2(n8611), .IN3(n7737), .IN4(n8644), .IN5(
        n7739), .IN6(n8846), .Q(n8610) );
  AO222X1 U8984 ( .IN1(n7747), .IN2(n8862), .IN3(n7743), .IN4(n8851), .IN5(
        n7745), .IN6(n8847), .Q(n8846) );
  AO222X1 U8985 ( .IN1(n8863), .IN2(n7626), .IN3(n8647), .IN4(n8852), .IN5(
        n7643), .IN6(n8848), .Q(n8847) );
  AO222X1 U8986 ( .IN1(n8699), .IN2(n8864), .IN3(n8697), .IN4(n8853), .IN5(
        n8711), .IN6(n8849), .Q(n8848) );
  AO222X1 U8987 ( .IN1(n8538), .IN2(n8865), .IN3(n8536), .IN4(n8854), .IN5(
        n8525), .IN6(n8850), .Q(n8849) );
  AO222X1 U8988 ( .IN1(n8767), .IN2(n7288), .IN3(n8779), .IN4(n7287), .IN5(
        n8766), .IN6(n7289), .Q(n8850) );
  INVX0 U8989 ( .INP(n4465), .ZN(n7287) );
  NOR2X0 U8990 ( .IN1(n7605), .IN2(n8368), .QN(n7739) );
  INVX0 U8991 ( .INP(n8083), .ZN(n7605) );
  AO222X1 U8992 ( .IN1(n7745), .IN2(n8851), .IN3(n7747), .IN4(n8645), .IN5(
        n7743), .IN6(n8862), .Q(n8644) );
  AO222X1 U8993 ( .IN1(n7643), .IN2(n8852), .IN3(n8866), .IN4(n7626), .IN5(
        n8647), .IN6(n8863), .Q(n8851) );
  AO222X1 U8994 ( .IN1(n8711), .IN2(n8853), .IN3(n8699), .IN4(n8867), .IN5(
        n8697), .IN6(n8864), .Q(n8852) );
  AO222X1 U8995 ( .IN1(n8525), .IN2(n8854), .IN3(n8538), .IN4(n8868), .IN5(
        n8536), .IN6(n8865), .Q(n8853) );
  AO222X1 U8996 ( .IN1(n8767), .IN2(n7289), .IN3(n8779), .IN4(n7288), .IN5(
        n8766), .IN6(n7290), .Q(n8854) );
  INVX0 U8997 ( .INP(n4464), .ZN(n7288) );
  XNOR2X1 U8998 ( .IN1(n8368), .IN2(n8083), .Q(n7737) );
  AO222X1 U8999 ( .IN1(n7747), .IN2(n8612), .IN3(n7743), .IN4(n8645), .IN5(
        n7745), .IN6(n8862), .Q(n8611) );
  AO222X1 U9000 ( .IN1(n8869), .IN2(n7626), .IN3(n8647), .IN4(n8866), .IN5(
        n7643), .IN6(n8863), .Q(n8862) );
  AO222X1 U9001 ( .IN1(n8699), .IN2(n8870), .IN3(n8697), .IN4(n8867), .IN5(
        n8711), .IN6(n8864), .Q(n8863) );
  AO222X1 U9002 ( .IN1(n8538), .IN2(n8871), .IN3(n8536), .IN4(n8868), .IN5(
        n8525), .IN6(n8865), .Q(n8864) );
  AO222X1 U9003 ( .IN1(n8767), .IN2(n7290), .IN3(n8779), .IN4(n7289), .IN5(
        n8766), .IN6(n7291), .Q(n8865) );
  INVX0 U9004 ( .INP(n4463), .ZN(n7289) );
  NOR2X0 U9005 ( .IN1(n8211), .IN2(n8369), .QN(n7745) );
  INVX0 U9006 ( .INP(n8380), .ZN(n8369) );
  AO222X1 U9007 ( .IN1(n7643), .IN2(n8866), .IN3(n8646), .IN4(n7626), .IN5(
        n8647), .IN6(n8869), .Q(n8645) );
  AO222X1 U9008 ( .IN1(n8711), .IN2(n8867), .IN3(n8699), .IN4(n8872), .IN5(
        n8697), .IN6(n8870), .Q(n8866) );
  AO222X1 U9009 ( .IN1(n8525), .IN2(n8868), .IN3(n8538), .IN4(n8873), .IN5(
        n8536), .IN6(n8871), .Q(n8867) );
  AO222X1 U9010 ( .IN1(n8767), .IN2(n7291), .IN3(n8779), .IN4(n7290), .IN5(
        n8766), .IN6(n7292), .Q(n8868) );
  INVX0 U9011 ( .INP(n4462), .ZN(n7290) );
  XNOR2X1 U9012 ( .IN1(n8211), .IN2(n8380), .Q(n7743) );
  AO222X1 U9013 ( .IN1(n8568), .IN2(n7626), .IN3(n8647), .IN4(n8646), .IN5(
        n7643), .IN6(n8869), .Q(n8612) );
  AO222X1 U9014 ( .IN1(n8699), .IN2(n8874), .IN3(n8697), .IN4(n8872), .IN5(
        n8711), .IN6(n8870), .Q(n8869) );
  AO222X1 U9015 ( .IN1(n8538), .IN2(n8875), .IN3(n8536), .IN4(n8873), .IN5(
        n8525), .IN6(n8871), .Q(n8870) );
  AO222X1 U9016 ( .IN1(n8767), .IN2(n7292), .IN3(n8779), .IN4(n7291), .IN5(
        n8766), .IN6(n7293), .Q(n8871) );
  INVX0 U9017 ( .INP(n4461), .ZN(n7291) );
  AO222X1 U9018 ( .IN1(n8711), .IN2(n8872), .IN3(n8699), .IN4(n8535), .IN5(
        n8697), .IN6(n8874), .Q(n8646) );
  AO222X1 U9019 ( .IN1(n8525), .IN2(n8873), .IN3(n8538), .IN4(n8876), .IN5(
        n8536), .IN6(n8875), .Q(n8872) );
  AO222X1 U9020 ( .IN1(n8767), .IN2(n7293), .IN3(n8779), .IN4(n7292), .IN5(
        n8766), .IN6(n7294), .Q(n8873) );
  INVX0 U9021 ( .INP(n4460), .ZN(n7292) );
  INVX0 U9022 ( .INP(n7749), .ZN(n8647) );
  NAND2X0 U9023 ( .IN1(n7751), .IN2(n7753), .QN(n7749) );
  AO221X1 U9024 ( .IN1(\r1720/A[3] ), .IN2(n8680), .IN3(n8877), .IN4(n8878), 
        .IN5(n8879), .Q(n7751) );
  AO222X1 U9025 ( .IN1(n8699), .IN2(n8523), .IN3(n8697), .IN4(n8535), .IN5(
        n8711), .IN6(n8874), .Q(n8568) );
  AO222X1 U9026 ( .IN1(n8538), .IN2(n8880), .IN3(n8536), .IN4(n8876), .IN5(
        n8525), .IN6(n8875), .Q(n8874) );
  AO222X1 U9027 ( .IN1(n8767), .IN2(n7294), .IN3(n8779), .IN4(n7293), .IN5(
        n8766), .IN6(n7295), .Q(n8875) );
  INVX0 U9028 ( .INP(n4459), .ZN(n7293) );
  INVX0 U9029 ( .INP(n7757), .ZN(n8711) );
  NAND2X0 U9030 ( .IN1(n7649), .IN2(n7625), .QN(n7757) );
  AO222X1 U9031 ( .IN1(n8525), .IN2(n8876), .IN3(n8538), .IN4(n8537), .IN5(
        n8536), .IN6(n8880), .Q(n8535) );
  AO222X1 U9032 ( .IN1(n8767), .IN2(n7295), .IN3(n8779), .IN4(n7294), .IN5(
        n8766), .IN6(n7296), .Q(n8876) );
  INVX0 U9033 ( .INP(n4458), .ZN(n7294) );
  XOR2X1 U9034 ( .IN1(n7649), .IN2(n7625), .Q(n8697) );
  AO222X1 U9035 ( .IN1(n8538), .IN2(n8524), .IN3(n8536), .IN4(n8537), .IN5(
        n8525), .IN6(n8880), .Q(n8523) );
  AO222X1 U9036 ( .IN1(n8767), .IN2(n7296), .IN3(n8779), .IN4(n7295), .IN5(
        n8766), .IN6(n7297), .Q(n8880) );
  INVX0 U9037 ( .INP(n4457), .ZN(n7295) );
  NOR2X0 U9038 ( .IN1(n8411), .IN2(n7660), .QN(n8525) );
  AO222X1 U9039 ( .IN1(n8767), .IN2(n7297), .IN3(n8779), .IN4(n7296), .IN5(
        n8766), .IN6(n7298), .Q(n8537) );
  INVX0 U9040 ( .INP(n7766), .ZN(n8766) );
  NAND2X0 U9041 ( .IN1(n8412), .IN2(n7666), .QN(n7766) );
  INVX0 U9042 ( .INP(n4456), .ZN(n7296) );
  INVX0 U9043 ( .INP(n7765), .ZN(n8767) );
  XOR2X1 U9044 ( .IN1(n8412), .IN2(n8078), .Q(n7765) );
  INVX0 U9045 ( .INP(n7666), .ZN(n8078) );
  INVX0 U9046 ( .INP(n7761), .ZN(n8536) );
  XNOR2X1 U9047 ( .IN1(n8411), .IN2(n7660), .Q(n7761) );
  MUX21X1 U9048 ( .IN1(n7298), .IN2(n7297), .S(n8779), .Q(n8524) );
  NOR2X0 U9049 ( .IN1(n7666), .IN2(n8412), .QN(n8779) );
  NAND3X0 U9050 ( .IN1(n8881), .IN2(n8882), .IN3(n8883), .QN(n8412) );
  NAND2X0 U9051 ( .IN1(\r1720/A[3] ), .IN2(n8884), .QN(n8882) );
  NAND3X0 U9052 ( .IN1(n8885), .IN2(n8886), .IN3(n8883), .QN(n7666) );
  NAND2X0 U9053 ( .IN1(\r1720/A[3] ), .IN2(n8887), .QN(n8885) );
  INVX0 U9054 ( .INP(n4455), .ZN(n7297) );
  INVX0 U9055 ( .INP(n4454), .ZN(n7298) );
  INVX0 U9056 ( .INP(n7764), .ZN(n8538) );
  NAND2X0 U9057 ( .IN1(n8411), .IN2(n7660), .QN(n7764) );
  NAND3X0 U9058 ( .IN1(n8888), .IN2(n8889), .IN3(n8890), .QN(n7660) );
  NAND2X0 U9059 ( .IN1(\r1720/A[3] ), .IN2(n8878), .QN(n8889) );
  NAND3X0 U9060 ( .IN1(n8881), .IN2(n8891), .IN3(n8883), .QN(n8411) );
  NOR2X0 U9061 ( .IN1(n8879), .IN2(n8877), .QN(n8883) );
  NAND3X0 U9062 ( .IN1(n8892), .IN2(n7526), .IN3(n8884), .QN(n8891) );
  INVX0 U9063 ( .INP(n8893), .ZN(n8884) );
  NOR2X0 U9064 ( .IN1(n7649), .IN2(n7625), .QN(n8699) );
  OA221X1 U9065 ( .IN1(n8886), .IN2(n7526), .IN3(n8894), .IN4(n8895), .IN5(
        n7753), .Q(n7625) );
  INVX0 U9066 ( .INP(n7626), .ZN(n7753) );
  OA221X1 U9067 ( .IN1(n7526), .IN2(n8890), .IN3(n8898), .IN4(n8899), .IN5(
        n8888), .Q(n7649) );
  NOR2X0 U9068 ( .IN1(n8877), .IN2(n8859), .QN(n8890) );
  NOR2X0 U9069 ( .IN1(n8225), .IN2(n8380), .QN(n7747) );
  OA21X1 U9070 ( .IN1(n8897), .IN2(n8899), .IN3(n8888), .Q(n8380) );
  INVX0 U9071 ( .INP(n8211), .ZN(n8225) );
  NAND4X0 U9072 ( .IN1(n8888), .IN2(n8900), .IN3(n8901), .IN4(n8902), .QN(
        n8211) );
  NAND2X0 U9073 ( .IN1(n8887), .IN2(n7526), .QN(n8901) );
  NAND2X0 U9074 ( .IN1(n8877), .IN2(n8718), .QN(n8900) );
  NOR2X0 U9075 ( .IN1(n8083), .IN2(n8381), .QN(n7741) );
  INVX0 U9076 ( .INP(n8368), .ZN(n8381) );
  NAND3X0 U9077 ( .IN1(n8903), .IN2(n8904), .IN3(n8888), .QN(n8368) );
  INVX0 U9078 ( .INP(n8879), .ZN(n8888) );
  NAND2X0 U9079 ( .IN1(n8855), .IN2(n8860), .QN(n8903) );
  INVX0 U9080 ( .INP(n8897), .ZN(n8855) );
  OA221X1 U9081 ( .IN1(n8897), .IN2(n8905), .IN3(n8906), .IN4(n8899), .IN5(
        n8861), .Q(n8083) );
  NAND2X0 U9082 ( .IN1(\r1720/A[3] ), .IN2(n8877), .QN(n8897) );
  AND2X1 U9083 ( .IN1(n8053), .IN2(n7650), .Q(n7733) );
  AO21X1 U9084 ( .IN1(n8907), .IN2(n8718), .IN3(n8879), .Q(n7650) );
  NAND2X0 U9085 ( .IN1(n8895), .IN2(n8908), .QN(n8879) );
  OAI21X1 U9086 ( .IN1(n8904), .IN2(n7526), .IN3(n8861), .QN(n8053) );
  NOR2X0 U9087 ( .IN1(n8683), .IN2(n8909), .QN(n8861) );
  NAND2X0 U9088 ( .IN1(n8678), .IN2(n8877), .QN(n8904) );
  AND2X1 U9089 ( .IN1(n8318), .IN2(n7644), .Q(n7724) );
  NAND3X0 U9090 ( .IN1(n8910), .IN2(n8911), .IN3(n8896), .QN(n7644) );
  AOI21X1 U9091 ( .IN1(n8857), .IN2(n8718), .IN3(n8679), .QN(n8896) );
  NAND2X0 U9092 ( .IN1(n8907), .IN2(n8860), .QN(n8911) );
  AO21X1 U9093 ( .IN1(n8909), .IN2(n8887), .IN3(n8912), .Q(n8318) );
  INVX0 U9094 ( .INP(n8899), .ZN(n8887) );
  NOR2X0 U9095 ( .IN1(n8913), .IN2(n8860), .QN(n8899) );
  AND2X1 U9096 ( .IN1(n8391), .IN2(n7671), .Q(n7718) );
  NAND4X0 U9097 ( .IN1(n8902), .IN2(n8906), .IN3(n8914), .IN4(n8915), .QN(
        n7671) );
  OA21X1 U9098 ( .IN1(n8895), .IN2(n8881), .IN3(n8910), .Q(n8915) );
  NAND2X0 U9099 ( .IN1(n8718), .IN2(n7526), .QN(n8914) );
  AO221X1 U9100 ( .IN1(n8916), .IN2(n8907), .IN3(n8857), .IN4(n8878), .IN5(
        n7638), .Q(n8391) );
  NOR2X0 U9101 ( .IN1(n8894), .IN2(n8881), .QN(n8916) );
  NOR2X0 U9102 ( .IN1(n8806), .IN2(n7706), .QN(n7709) );
  NOR2X0 U9103 ( .IN1(n8912), .IN2(n8917), .QN(n7706) );
  AND3X1 U9104 ( .IN1(n8860), .IN2(n8892), .IN3(n8918), .Q(n8917) );
  NAND3X0 U9105 ( .IN1(n8906), .IN2(n8908), .IN3(n8919), .QN(n8912) );
  NAND2X0 U9106 ( .IN1(n8859), .IN2(n8857), .QN(n8919) );
  INVX0 U9107 ( .INP(n7712), .ZN(n8806) );
  AO221X1 U9108 ( .IN1(n8909), .IN2(n8856), .IN3(n8679), .IN4(\r1720/A[3] ), 
        .IN5(n8719), .Q(n7712) );
  AO21X1 U9109 ( .IN1(n8859), .IN2(n8679), .IN3(n8683), .Q(n8719) );
  AND2X1 U9110 ( .IN1(n8227), .IN2(n7638), .Q(n7701) );
  NAND3X0 U9111 ( .IN1(n8920), .IN2(n8906), .IN3(n8910), .QN(n7638) );
  NAND2X0 U9112 ( .IN1(n8859), .IN2(n8907), .QN(n8920) );
  INVX0 U9113 ( .INP(n8902), .ZN(n8907) );
  NAND3X0 U9114 ( .IN1(n8717), .IN2(n8908), .IN3(n8921), .QN(n8227) );
  NAND2X0 U9115 ( .IN1(n8909), .IN2(n8680), .QN(n8921) );
  OR2X1 U9116 ( .IN1(n8877), .IN2(n8678), .Q(n8680) );
  AND2X1 U9117 ( .IN1(n8859), .IN2(n8892), .Q(n8678) );
  INVX0 U9118 ( .INP(n8894), .ZN(n8892) );
  NOR2X0 U9119 ( .IN1(n8881), .IN2(n8893), .QN(n8859) );
  NOR2X0 U9120 ( .IN1(n7526), .IN2(n8895), .QN(n8909) );
  NAND2X0 U9121 ( .IN1(n8856), .IN2(n8679), .QN(n8717) );
  INVX0 U9122 ( .INP(n8886), .ZN(n8856) );
  NAND2X0 U9123 ( .IN1(n8860), .IN2(n8913), .QN(n8886) );
  NOR2X0 U9124 ( .IN1(n8768), .IN2(n8353), .QN(n7694) );
  INVX0 U9125 ( .INP(n8337), .ZN(n8353) );
  AO221X1 U9126 ( .IN1(n8918), .IN2(n8860), .IN3(n8679), .IN4(n8718), .IN5(
        n8922), .Q(n8337) );
  NAND2X0 U9127 ( .IN1(n8893), .IN2(n8881), .QN(n8718) );
  INVX0 U9128 ( .INP(n8923), .ZN(n8918) );
  AO21X1 U9129 ( .IN1(n8905), .IN2(n8924), .IN3(n8906), .Q(n8768) );
  NAND2X0 U9130 ( .IN1(\r1720/A[3] ), .IN2(n8913), .QN(n8924) );
  NAND2X0 U9131 ( .IN1(n8894), .IN2(n8893), .QN(n8913) );
  NOR2X0 U9132 ( .IN1(n7692), .IN2(n8409), .QN(n7688) );
  INVX0 U9133 ( .INP(n8406), .ZN(n8409) );
  NAND3X0 U9134 ( .IN1(n8925), .IN2(n8902), .IN3(n8910), .QN(n8406) );
  INVX0 U9135 ( .INP(n8681), .ZN(n8910) );
  NAND2X0 U9136 ( .IN1(n8908), .IN2(n8923), .QN(n8681) );
  NAND2X0 U9137 ( .IN1(n8877), .IN2(n7526), .QN(n8902) );
  NAND2X0 U9138 ( .IN1(n8679), .IN2(n8860), .QN(n8925) );
  INVX0 U9139 ( .INP(n8881), .ZN(n8860) );
  INVX0 U9140 ( .INP(n8906), .ZN(n8679) );
  INVX0 U9141 ( .INP(n8338), .ZN(n7692) );
  AO21X1 U9142 ( .IN1(n8926), .IN2(n8878), .IN3(n8922), .Q(n8338) );
  INVX0 U9143 ( .INP(n8716), .ZN(n8922) );
  NOR2X0 U9144 ( .IN1(n8683), .IN2(n8682), .QN(n8716) );
  NOR2X0 U9145 ( .IN1(n8906), .IN2(\r1720/A[3] ), .QN(n8682) );
  INVX0 U9146 ( .INP(n8908), .ZN(n8683) );
  NAND2X0 U9147 ( .IN1(n8049), .IN2(n7526), .QN(n8908) );
  NAND3X0 U9148 ( .IN1(n4479), .IN2(n4478), .IN3(n4480), .QN(n8049) );
  INVX0 U9149 ( .INP(n8905), .ZN(n8878) );
  OA21X1 U9150 ( .IN1(n8893), .IN2(n8894), .IN3(n8881), .Q(n8905) );
  MUX21X1 U9151 ( .IN1(n4483), .IN2(n3715), .S(\r1720/A[3] ), .Q(n8881) );
  MUX21X1 U9152 ( .IN1(n4485), .IN2(n3713), .S(\r1720/A[3] ), .Q(n8894) );
  MUX21X1 U9153 ( .IN1(n4484), .IN2(n3714), .S(\r1720/A[3] ), .Q(n8893) );
  NAND2X0 U9154 ( .IN1(n8906), .IN2(n8923), .QN(n8926) );
  NAND2X0 U9155 ( .IN1(n8857), .IN2(n7526), .QN(n8923) );
  INVX0 U9156 ( .INP(\r1720/A[3] ), .ZN(n7526) );
  NAND2X0 U9157 ( .IN1(n8857), .IN2(n8877), .QN(n8906) );
  INVX0 U9158 ( .INP(n8898), .ZN(n8877) );
  MUX21X1 U9159 ( .IN1(n4482), .IN2(n3627), .S(\r1720/A[3] ), .Q(n8898) );
  INVX0 U9160 ( .INP(n8895), .ZN(n8857) );
  MUX21X1 U9161 ( .IN1(n4481), .IN2(n3628), .S(\r1720/A[3] ), .Q(n8895) );
  NOR2X0 U9162 ( .IN1(n4485), .IN2(n3630), .QN(N1895) );
  NOR2X0 U9163 ( .IN1(n4484), .IN2(n3631), .QN(N1894) );
  NOR2X0 U9164 ( .IN1(n4483), .IN2(n3632), .QN(N1893) );
  NOR2X0 U9165 ( .IN1(n4482), .IN2(n3633), .QN(N1892) );
  NOR2X0 U9166 ( .IN1(n4481), .IN2(n3634), .QN(N1891) );
  NOR2X0 U9167 ( .IN1(n4480), .IN2(n3635), .QN(N1890) );
  NOR2X0 U9168 ( .IN1(n4479), .IN2(n3636), .QN(N1889) );
  NOR2X0 U9169 ( .IN1(n4478), .IN2(n3637), .QN(N1888) );
  NOR2X0 U9170 ( .IN1(n4477), .IN2(n3638), .QN(N1887) );
  NOR2X0 U9171 ( .IN1(n4476), .IN2(n3639), .QN(N1886) );
  NOR2X0 U9172 ( .IN1(n4475), .IN2(n3640), .QN(N1885) );
  NOR2X0 U9173 ( .IN1(n4474), .IN2(n3641), .QN(N1884) );
  NOR2X0 U9174 ( .IN1(n4473), .IN2(n3642), .QN(N1883) );
  NOR2X0 U9175 ( .IN1(n4472), .IN2(n3643), .QN(N1882) );
  NOR2X0 U9176 ( .IN1(n4471), .IN2(n3644), .QN(N1881) );
  NOR2X0 U9177 ( .IN1(n4470), .IN2(n3645), .QN(N1880) );
  NOR2X0 U9178 ( .IN1(n4469), .IN2(n3646), .QN(N1879) );
  NOR2X0 U9179 ( .IN1(n4468), .IN2(n3647), .QN(N1878) );
  NOR2X0 U9180 ( .IN1(n4467), .IN2(n3648), .QN(N1877) );
  NOR2X0 U9181 ( .IN1(n4466), .IN2(n3649), .QN(N1876) );
  NOR2X0 U9182 ( .IN1(n4465), .IN2(n3650), .QN(N1875) );
  NOR2X0 U9183 ( .IN1(n4464), .IN2(n3651), .QN(N1874) );
  NOR2X0 U9184 ( .IN1(n4463), .IN2(n3652), .QN(N1873) );
  NOR2X0 U9185 ( .IN1(n4462), .IN2(n3653), .QN(N1872) );
  NOR2X0 U9186 ( .IN1(n4461), .IN2(n3654), .QN(N1871) );
  NOR2X0 U9187 ( .IN1(n4460), .IN2(n3655), .QN(N1870) );
  NOR2X0 U9188 ( .IN1(n4459), .IN2(n3656), .QN(N1869) );
  NOR2X0 U9189 ( .IN1(n4458), .IN2(n3657), .QN(N1868) );
  NOR2X0 U9190 ( .IN1(n4457), .IN2(n3658), .QN(N1867) );
  NOR2X0 U9191 ( .IN1(n4456), .IN2(n3659), .QN(N1866) );
  NOR2X0 U9192 ( .IN1(n4455), .IN2(n3660), .QN(N1865) );
  NOR2X0 U9193 ( .IN1(n4454), .IN2(n3661), .QN(N1864) );
  NOR2X0 U9194 ( .IN1(n3693), .IN2(n4485), .QN(N1255) );
  NOR2X0 U9195 ( .IN1(n3692), .IN2(n4484), .QN(N1254) );
  NAND4X0 U9196 ( .IN1(n8927), .IN2(n8928), .IN3(n8929), .IN4(n8930), .QN(
        N1192) );
  NOR4X0 U9197 ( .IN1(n8931), .IN2(n8932), .IN3(n8933), .IN4(n8934), .QN(n8930) );
  INVX0 U9198 ( .INP(n8935), .ZN(n8934) );
  AO22X1 U9199 ( .IN1(n7346), .IN2(n5702), .IN3(n7308), .IN4(n8936), .Q(n8931)
         );
  NAND4X0 U9200 ( .IN1(n8937), .IN2(n7312), .IN3(n7368), .IN4(n8938), .QN(
        n8936) );
  NOR2X0 U9201 ( .IN1(n8939), .IN2(n8940), .QN(n8938) );
  AOI21X1 U9202 ( .IN1(n7355), .IN2(n7363), .IN3(n7362), .QN(n8939) );
  NAND2X0 U9203 ( .IN1(n7223), .IN2(n8941), .QN(n7346) );
  OA222X1 U9204 ( .IN1(n7364), .IN2(n7350), .IN3(n8942), .IN4(n7348), .IN5(
        n3711), .IN6(n7300), .Q(n8929) );
  NAND4X0 U9205 ( .IN1(n8943), .IN2(n8944), .IN3(n8945), .IN4(n8946), .QN(
        N1191) );
  OA221X1 U9206 ( .IN1(n7123), .IN2(n8947), .IN3(n5702), .IN4(n7348), .IN5(
        n8948), .Q(n8946) );
  OA21X1 U9207 ( .IN1(n8949), .IN2(n7223), .IN3(n8950), .Q(n8948) );
  NOR3X0 U9208 ( .IN1(n7373), .IN2(n8933), .IN3(n8951), .QN(n8945) );
  AND3X1 U9209 ( .IN1(n8952), .IN2(n8953), .IN3(n7340), .Q(n8951) );
  NAND3X0 U9210 ( .IN1(n4422), .IN2(n7129), .IN3(n8954), .QN(n8944) );
  NAND2X0 U9211 ( .IN1(n7308), .IN2(n8955), .QN(n8943) );
  NAND4X0 U9212 ( .IN1(n8956), .IN2(n7367), .IN3(n4422), .IN4(n7310), .QN(
        n8955) );
  INVX0 U9213 ( .INP(n8957), .ZN(n7367) );
  INVX0 U9214 ( .INP(n8958), .ZN(n8956) );
  NAND4X0 U9215 ( .IN1(n8927), .IN2(n8959), .IN3(n8960), .IN4(n8961), .QN(
        N1190) );
  OA221X1 U9216 ( .IN1(n9186), .IN2(n7350), .IN3(n8962), .IN4(n7142), .IN5(
        n8963), .Q(n8961) );
  NOR2X0 U9217 ( .IN1(n8964), .IN2(n8965), .QN(n8963) );
  AOI21X1 U9218 ( .IN1(n8966), .IN2(n7123), .IN3(n8947), .QN(n8965) );
  INVX0 U9219 ( .INP(n8932), .ZN(n8947) );
  NOR4X0 U9220 ( .IN1(n8967), .IN2(n8968), .IN3(n8940), .IN4(n8958), .QN(n8962) );
  NAND3X0 U9221 ( .IN1(n7370), .IN2(n7147), .IN3(n7356), .QN(n8958) );
  AO22X1 U9222 ( .IN1(n8969), .IN2(n8970), .IN3(n8971), .IN4(n8972), .Q(n8968)
         );
  NAND4X0 U9223 ( .IN1(n8973), .IN2(n7312), .IN3(n7311), .IN4(n7343), .QN(
        n8967) );
  MUX21X1 U9224 ( .IN1(n8974), .IN2(n8941), .S(n7226), .Q(n8960) );
  NAND2X0 U9225 ( .IN1(n8975), .IN2(n8953), .QN(n8959) );
  AOI21X1 U9226 ( .IN1(n8954), .IN2(n8976), .IN3(n9191), .QN(n8927) );
  OR3X1 U9227 ( .IN1(n7107), .IN2(n7345), .IN3(n7129), .Q(n8976) );
  NAND4X0 U9228 ( .IN1(n7344), .IN2(n8977), .IN3(n8978), .IN4(n8979), .QN(
        N1189) );
  NOR4X0 U9229 ( .IN1(n8980), .IN2(n8981), .IN3(n8982), .IN4(n8983), .QN(n8979) );
  MUX21X1 U9230 ( .IN1(n8975), .IN2(n8964), .S(n9187), .Q(n8983) );
  INVX0 U9231 ( .INP(n8928), .ZN(n8980) );
  OA21X1 U9232 ( .IN1(n8974), .IN2(n8984), .IN3(n8985), .Q(n8928) );
  NAND4X0 U9233 ( .IN1(n8971), .IN2(n7308), .IN3(n7129), .IN4(n7105), .QN(
        n8985) );
  INVX0 U9234 ( .INP(n7355), .ZN(n8971) );
  OA221X1 U9235 ( .IN1(n8986), .IN2(n7142), .IN3(n8987), .IN4(n7307), .IN5(
        n8988), .Q(n8978) );
  NAND3X0 U9236 ( .IN1(n8952), .IN2(n8953), .IN3(n7306), .QN(n8988) );
  NAND2X0 U9237 ( .IN1(n3711), .IN2(n8984), .QN(n8952) );
  NOR2X0 U9238 ( .IN1(n7222), .IN2(n7373), .QN(n8987) );
  INVX0 U9239 ( .INP(n7348), .ZN(n7222) );
  OA221X1 U9240 ( .IN1(n7363), .IN2(n8970), .IN3(n3697), .IN4(n7361), .IN5(
        n8989), .Q(n8986) );
  NOR2X0 U9241 ( .IN1(n8957), .IN2(n8990), .QN(n8989) );
  NAND4X0 U9242 ( .IN1(n8937), .IN2(n8973), .IN3(n8991), .IN4(n7343), .QN(
        n8957) );
  NAND2X0 U9243 ( .IN1(n8992), .IN2(n7126), .QN(n8973) );
  NAND3X0 U9244 ( .IN1(n4422), .IN2(n7105), .IN3(n8992), .QN(n8937) );
  NOR2X0 U9245 ( .IN1(n8969), .IN2(n8993), .QN(n7363) );
  INVX0 U9246 ( .INP(n7361), .ZN(n8969) );
  NAND2X0 U9247 ( .IN1(n8933), .IN2(n3700), .QN(n8977) );
  OA21X1 U9248 ( .IN1(n7140), .IN2(n9187), .IN3(n7143), .Q(n7344) );
  NAND4X0 U9249 ( .IN1(n8994), .IN2(n8950), .IN3(n8995), .IN4(n8996), .QN(
        N1188) );
  OA221X1 U9250 ( .IN1(n7107), .IN2(n7300), .IN3(n7226), .IN4(n7348), .IN5(
        n8997), .Q(n8996) );
  OA222X1 U9251 ( .IN1(n8998), .IN2(n7142), .IN3(n8999), .IN4(n7117), .IN5(
        n9000), .IN6(n8984), .Q(n8997) );
  NOR2X0 U9252 ( .IN1(n7306), .IN2(n8975), .QN(n9000) );
  INVX0 U9253 ( .INP(n7223), .ZN(n8975) );
  NOR2X0 U9254 ( .IN1(n3700), .IN2(n7128), .QN(n8999) );
  OA21X1 U9255 ( .IN1(n8970), .IN2(n7361), .IN3(n9001), .Q(n8998) );
  NAND2X0 U9256 ( .IN1(n7227), .IN2(n5692), .QN(n7348) );
  OA222X1 U9257 ( .IN1(n3700), .IN2(n7145), .IN3(n8942), .IN4(n7342), .IN5(
        n8992), .IN6(n8941), .Q(n8995) );
  INVX0 U9258 ( .INP(n8953), .ZN(n8942) );
  AND4X1 U9259 ( .IN1(n9002), .IN2(n9003), .IN3(n9004), .IN4(n7143), .Q(n8950)
         );
  NAND2X0 U9260 ( .IN1(n7226), .IN2(n7308), .QN(n7143) );
  NAND2X0 U9261 ( .IN1(n7308), .IN2(n9005), .QN(n9004) );
  NAND3X0 U9262 ( .IN1(n7368), .IN2(n7312), .IN3(n9006), .QN(n9005) );
  NAND2X0 U9263 ( .IN1(n9007), .IN2(n8993), .QN(n9006) );
  NAND2X0 U9264 ( .IN1(n9008), .IN2(n9009), .QN(n7312) );
  NAND2X0 U9265 ( .IN1(n8992), .IN2(n7123), .QN(n7368) );
  INVX0 U9266 ( .INP(n9010), .ZN(n8992) );
  NAND2X0 U9267 ( .IN1(n7226), .IN2(n7221), .QN(n9003) );
  INVX0 U9268 ( .INP(n8982), .ZN(n8994) );
  AO22X1 U9269 ( .IN1(n8932), .IN2(n8966), .IN3(n9011), .IN4(n3697), .Q(n8982)
         );
  NOR2X0 U9270 ( .IN1(n7107), .IN2(n7145), .QN(n9011) );
  NAND4X0 U9271 ( .IN1(n9002), .IN2(n9012), .IN3(n9013), .IN4(n9014), .QN(
        N1187) );
  NOR4X0 U9272 ( .IN1(n9015), .IN2(n9016), .IN3(n8933), .IN4(n7337), .QN(n9014) );
  INVX0 U9273 ( .INP(n7300), .ZN(n7337) );
  NAND2X0 U9274 ( .IN1(n7306), .IN2(n9017), .QN(n7300) );
  INVX0 U9275 ( .INP(n7350), .ZN(n7306) );
  NAND2X0 U9276 ( .IN1(n7340), .IN2(n5705), .QN(n7350) );
  NOR2X0 U9277 ( .IN1(n7128), .IN2(n7117), .QN(n8933) );
  NAND2X0 U9278 ( .IN1(n7221), .IN2(n9187), .QN(n7117) );
  INVX0 U9279 ( .INP(n8974), .ZN(n7221) );
  NAND2X0 U9280 ( .IN1(n7126), .IN2(n9186), .QN(n7128) );
  NOR3X0 U9281 ( .IN1(n7145), .IN2(n4422), .IN3(n7026), .QN(n9016) );
  INVX0 U9282 ( .INP(n8954), .ZN(n7145) );
  AO222X1 U9283 ( .IN1(n7373), .IN2(n8953), .IN3(n8932), .IN4(n8966), .IN5(
        n7308), .IN6(n9018), .Q(n9015) );
  NAND4X0 U9284 ( .IN1(n8991), .IN2(n7310), .IN3(n9019), .IN4(n9020), .QN(
        n9018) );
  OA221X1 U9285 ( .IN1(n7362), .IN2(n9021), .IN3(n7360), .IN4(n7361), .IN5(
        n9001), .Q(n9020) );
  AND3X1 U9286 ( .IN1(n9022), .IN2(n7370), .IN3(n9023), .Q(n9001) );
  INVX0 U9287 ( .INP(n8990), .ZN(n9023) );
  NAND4X0 U9288 ( .IN1(n9024), .IN2(n9025), .IN3(n7356), .IN4(n7311), .QN(
        n8990) );
  NAND3X0 U9289 ( .IN1(n7129), .IN2(n7105), .IN3(n8993), .QN(n7311) );
  INVX0 U9290 ( .INP(n9021), .ZN(n8993) );
  NAND2X0 U9291 ( .IN1(n8972), .IN2(n9009), .QN(n7356) );
  NAND2X0 U9292 ( .IN1(n9007), .IN2(n9009), .QN(n9025) );
  INVX0 U9293 ( .INP(n7360), .ZN(n9007) );
  INVX0 U9294 ( .INP(n8940), .ZN(n9024) );
  AO21X1 U9295 ( .IN1(n8949), .IN2(n7107), .IN3(n7372), .Q(n8940) );
  NOR3X0 U9296 ( .IN1(n7105), .IN2(n7107), .IN3(n9010), .QN(n7372) );
  NAND3X0 U9297 ( .IN1(n4422), .IN2(n7105), .IN3(n9017), .QN(n7370) );
  OR2X1 U9298 ( .IN1(n7355), .IN2(n7362), .Q(n9022) );
  NAND2X0 U9299 ( .IN1(n9026), .IN2(n6950), .QN(n7355) );
  NAND2X0 U9300 ( .IN1(n9026), .IN2(n3695), .QN(n7361) );
  NOR3X0 U9301 ( .IN1(n7107), .IN2(n3700), .IN3(n8984), .QN(n9026) );
  NAND2X0 U9302 ( .IN1(n3697), .IN2(n3711), .QN(n7360) );
  NAND4X0 U9303 ( .IN1(n8949), .IN2(n3700), .IN3(n4422), .IN4(n6946), .QN(
        n9021) );
  NOR2X0 U9304 ( .IN1(n9008), .IN2(n8972), .QN(n7362) );
  NOR2X0 U9305 ( .IN1(n7105), .IN2(n3697), .QN(n8972) );
  INVX0 U9306 ( .INP(n8970), .ZN(n9008) );
  NAND2X0 U9307 ( .IN1(n3697), .IN2(n7105), .QN(n8970) );
  AND2X1 U9308 ( .IN1(n7343), .IN2(n7147), .Q(n9019) );
  NAND2X0 U9309 ( .IN1(n7123), .IN2(n9017), .QN(n7147) );
  NAND2X0 U9310 ( .IN1(n9017), .IN2(n7126), .QN(n7343) );
  NOR2X0 U9311 ( .IN1(n4422), .IN2(n3711), .QN(n7126) );
  NAND3X0 U9312 ( .IN1(n7129), .IN2(n7105), .IN3(n9009), .QN(n7310) );
  INVX0 U9313 ( .INP(n7359), .ZN(n9009) );
  NAND4X0 U9314 ( .IN1(n3695), .IN2(n8949), .IN3(n3700), .IN4(n4422), .QN(
        n7359) );
  INVX0 U9315 ( .INP(n8984), .ZN(n8949) );
  INVX0 U9316 ( .INP(n3697), .ZN(n7129) );
  NAND3X0 U9317 ( .IN1(n3711), .IN2(n4422), .IN3(n9017), .QN(n8991) );
  INVX0 U9318 ( .INP(n7307), .ZN(n9017) );
  INVX0 U9319 ( .INP(n7142), .ZN(n7308) );
  NAND3X0 U9320 ( .IN1(n5686), .IN2(n5705), .IN3(n9188), .QN(n7142) );
  NAND2X0 U9321 ( .IN1(n7123), .IN2(n7016), .QN(n8966) );
  INVX0 U9322 ( .INP(n7146), .ZN(n7123) );
  NOR2X0 U9323 ( .IN1(n7140), .IN2(n7307), .QN(n8932) );
  NAND2X0 U9324 ( .IN1(n7307), .IN2(n8984), .QN(n8953) );
  NAND2X0 U9325 ( .IN1(n5702), .IN2(n5689), .QN(n8984) );
  NAND2X0 U9326 ( .IN1(n9187), .IN2(n9186), .QN(n7307) );
  INVX0 U9327 ( .INP(n8941), .ZN(n7373) );
  NAND2X0 U9328 ( .IN1(n7340), .IN2(n9185), .QN(n8941) );
  INVX0 U9329 ( .INP(n7365), .ZN(n7340) );
  NAND2X0 U9330 ( .IN1(n5692), .IN2(n5686), .QN(n7365) );
  OA222X1 U9331 ( .IN1(n7364), .IN2(n7140), .IN3(n9187), .IN4(n8974), .IN5(
        n9010), .IN6(n7223), .Q(n9013) );
  NAND2X0 U9332 ( .IN1(n7227), .IN2(n9188), .QN(n7223) );
  INVX0 U9333 ( .INP(n7141), .ZN(n7227) );
  NAND2X0 U9334 ( .IN1(n9189), .IN2(n5705), .QN(n7141) );
  NAND3X0 U9335 ( .IN1(n9188), .IN2(n5686), .IN3(n9185), .QN(n8974) );
  NAND2X0 U9336 ( .IN1(n8964), .IN2(n5702), .QN(n9012) );
  INVX0 U9337 ( .INP(n8981), .ZN(n9002) );
  NAND3X0 U9338 ( .IN1(n8935), .IN2(n5701), .IN3(n9027), .QN(n8981) );
  NAND2X0 U9339 ( .IN1(n7345), .IN2(n8954), .QN(n9027) );
  NOR2X0 U9340 ( .IN1(n9010), .IN2(n7140), .QN(n8954) );
  NAND3X0 U9341 ( .IN1(n9185), .IN2(n5692), .IN3(n9189), .QN(n7140) );
  NAND2X0 U9342 ( .IN1(n9187), .IN2(n5702), .QN(n9010) );
  OA21X1 U9343 ( .IN1(n7026), .IN2(n7105), .IN3(n7146), .Q(n7345) );
  NAND2X0 U9344 ( .IN1(n3711), .IN2(n7107), .QN(n7146) );
  INVX0 U9345 ( .INP(n4422), .ZN(n7107) );
  INVX0 U9346 ( .INP(n3711), .ZN(n7105) );
  NAND2X0 U9347 ( .IN1(n7226), .IN2(n8964), .QN(n8935) );
  INVX0 U9348 ( .INP(n7342), .ZN(n8964) );
  NAND3X0 U9349 ( .IN1(n9185), .IN2(n9188), .IN3(n9189), .QN(n7342) );
  INVX0 U9350 ( .INP(n7364), .ZN(n7226) );
  NAND2X0 U9351 ( .IN1(n9186), .IN2(n5689), .QN(n7364) );
endmodule



module pipealu_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [33:0] carry;
  wire   [32:0] B_AS;
  assign carry[0] = ADD_SUB;

  FADDX1 U1_31 ( .A(A[31]), .B(B_AS[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B_AS[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B_AS[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B_AS[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B_AS[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B_AS[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B_AS[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B_AS[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B_AS[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B_AS[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B_AS[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B_AS[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B_AS[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B_AS[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B_AS[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B_AS[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B_AS[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FADDX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FADDX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FADDX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FADDX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FADDX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FADDX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FADDX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FADDX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0]) );
  XOR2X1 U1 ( .IN1(carry[0]), .IN2(carry[32]), .Q(SUM[32]) );
  XOR2X1 U2 ( .IN1(B[9]), .IN2(carry[0]), .Q(B_AS[9]) );
  XOR2X1 U3 ( .IN1(B[8]), .IN2(carry[0]), .Q(B_AS[8]) );
  XOR2X1 U4 ( .IN1(B[7]), .IN2(carry[0]), .Q(B_AS[7]) );
  XOR2X1 U5 ( .IN1(B[6]), .IN2(carry[0]), .Q(B_AS[6]) );
  XOR2X1 U6 ( .IN1(B[5]), .IN2(carry[0]), .Q(B_AS[5]) );
  XOR2X1 U7 ( .IN1(B[4]), .IN2(carry[0]), .Q(B_AS[4]) );
  XOR2X1 U8 ( .IN1(B[3]), .IN2(carry[0]), .Q(B_AS[3]) );
  XOR2X1 U9 ( .IN1(B[31]), .IN2(carry[0]), .Q(B_AS[31]) );
  XOR2X1 U10 ( .IN1(B[30]), .IN2(carry[0]), .Q(B_AS[30]) );
  XOR2X1 U11 ( .IN1(B[2]), .IN2(carry[0]), .Q(B_AS[2]) );
  XOR2X1 U12 ( .IN1(B[29]), .IN2(carry[0]), .Q(B_AS[29]) );
  XOR2X1 U13 ( .IN1(B[28]), .IN2(carry[0]), .Q(B_AS[28]) );
  XOR2X1 U14 ( .IN1(B[27]), .IN2(carry[0]), .Q(B_AS[27]) );
  XOR2X1 U15 ( .IN1(B[26]), .IN2(carry[0]), .Q(B_AS[26]) );
  XOR2X1 U16 ( .IN1(B[25]), .IN2(carry[0]), .Q(B_AS[25]) );
  XOR2X1 U17 ( .IN1(B[24]), .IN2(carry[0]), .Q(B_AS[24]) );
  XOR2X1 U18 ( .IN1(B[23]), .IN2(carry[0]), .Q(B_AS[23]) );
  XOR2X1 U19 ( .IN1(B[22]), .IN2(carry[0]), .Q(B_AS[22]) );
  XOR2X1 U20 ( .IN1(B[21]), .IN2(carry[0]), .Q(B_AS[21]) );
  XOR2X1 U21 ( .IN1(B[20]), .IN2(carry[0]), .Q(B_AS[20]) );
  XOR2X1 U22 ( .IN1(B[1]), .IN2(carry[0]), .Q(B_AS[1]) );
  XOR2X1 U23 ( .IN1(B[19]), .IN2(carry[0]), .Q(B_AS[19]) );
  XOR2X1 U24 ( .IN1(B[18]), .IN2(carry[0]), .Q(B_AS[18]) );
  XOR2X1 U25 ( .IN1(B[17]), .IN2(carry[0]), .Q(B_AS[17]) );
  XOR2X1 U26 ( .IN1(B[16]), .IN2(carry[0]), .Q(B_AS[16]) );
  XOR2X1 U27 ( .IN1(B[15]), .IN2(carry[0]), .Q(B_AS[15]) );
  XOR2X1 U28 ( .IN1(B[14]), .IN2(carry[0]), .Q(B_AS[14]) );
  XOR2X1 U29 ( .IN1(B[13]), .IN2(carry[0]), .Q(B_AS[13]) );
  XOR2X1 U30 ( .IN1(B[12]), .IN2(carry[0]), .Q(B_AS[12]) );
  XOR2X1 U31 ( .IN1(B[11]), .IN2(carry[0]), .Q(B_AS[11]) );
  XOR2X1 U32 ( .IN1(B[10]), .IN2(carry[0]), .Q(B_AS[10]) );
  XOR2X1 U33 ( .IN1(B[0]), .IN2(carry[0]), .Q(B_AS[0]) );
endmodule


module pipealu ( instr, AluOut, Zero, clk, Carryout, Overflow, rst );
  input [15:0] instr;
  output [31:0] AluOut;
  input clk, rst;
  output Zero, Carryout, Overflow;
  wire   N15, N16, N17, N18, N19, N20, N21, N22, \regfile[15][31] ,
         \regfile[15][30] , \regfile[15][29] , \regfile[15][28] ,
         \regfile[15][27] , \regfile[15][26] , \regfile[15][25] ,
         \regfile[15][24] , \regfile[15][23] , \regfile[15][22] ,
         \regfile[15][21] , \regfile[15][20] , \regfile[15][19] ,
         \regfile[15][18] , \regfile[15][17] , \regfile[15][16] ,
         \regfile[15][15] , \regfile[15][14] , \regfile[15][13] ,
         \regfile[15][12] , \regfile[15][11] , \regfile[15][10] ,
         \regfile[15][9] , \regfile[15][8] , \regfile[15][7] ,
         \regfile[15][6] , \regfile[15][5] , \regfile[15][4] ,
         \regfile[15][3] , \regfile[15][2] , \regfile[15][1] ,
         \regfile[15][0] , \regfile[14][31] , \regfile[14][30] ,
         \regfile[14][29] , \regfile[14][28] , \regfile[14][27] ,
         \regfile[14][26] , \regfile[14][25] , \regfile[14][24] ,
         \regfile[14][23] , \regfile[14][22] , \regfile[14][21] ,
         \regfile[14][20] , \regfile[14][19] , \regfile[14][18] ,
         \regfile[14][17] , \regfile[14][16] , \regfile[14][15] ,
         \regfile[14][14] , \regfile[14][13] , \regfile[14][12] ,
         \regfile[14][11] , \regfile[14][10] , \regfile[14][9] ,
         \regfile[14][8] , \regfile[14][7] , \regfile[14][6] ,
         \regfile[14][5] , \regfile[14][4] , \regfile[14][3] ,
         \regfile[14][2] , \regfile[14][1] , \regfile[14][0] ,
         \regfile[13][31] , \regfile[13][30] , \regfile[13][29] ,
         \regfile[13][28] , \regfile[13][27] , \regfile[13][26] ,
         \regfile[13][25] , \regfile[13][24] , \regfile[13][23] ,
         \regfile[13][22] , \regfile[13][21] , \regfile[13][20] ,
         \regfile[13][19] , \regfile[13][18] , \regfile[13][17] ,
         \regfile[13][16] , \regfile[13][15] , \regfile[13][14] ,
         \regfile[13][13] , \regfile[13][12] , \regfile[13][11] ,
         \regfile[13][10] , \regfile[13][9] , \regfile[13][8] ,
         \regfile[13][7] , \regfile[13][6] , \regfile[13][5] ,
         \regfile[13][4] , \regfile[13][3] , \regfile[13][2] ,
         \regfile[13][1] , \regfile[13][0] , \regfile[12][31] ,
         \regfile[12][30] , \regfile[12][29] , \regfile[12][28] ,
         \regfile[12][27] , \regfile[12][26] , \regfile[12][25] ,
         \regfile[12][24] , \regfile[12][23] , \regfile[12][22] ,
         \regfile[12][21] , \regfile[12][20] , \regfile[12][19] ,
         \regfile[12][18] , \regfile[12][17] , \regfile[12][16] ,
         \regfile[12][15] , \regfile[12][14] , \regfile[12][13] ,
         \regfile[12][12] , \regfile[12][11] , \regfile[12][10] ,
         \regfile[12][9] , \regfile[12][8] , \regfile[12][7] ,
         \regfile[12][6] , \regfile[12][5] , \regfile[12][4] ,
         \regfile[12][3] , \regfile[12][2] , \regfile[12][1] ,
         \regfile[12][0] , \regfile[11][31] , \regfile[11][30] ,
         \regfile[11][29] , \regfile[11][28] , \regfile[11][27] ,
         \regfile[11][26] , \regfile[11][25] , \regfile[11][24] ,
         \regfile[11][23] , \regfile[11][22] , \regfile[11][21] ,
         \regfile[11][20] , \regfile[11][19] , \regfile[11][18] ,
         \regfile[11][17] , \regfile[11][16] , \regfile[11][15] ,
         \regfile[11][14] , \regfile[11][13] , \regfile[11][12] ,
         \regfile[11][11] , \regfile[11][10] , \regfile[11][9] ,
         \regfile[11][8] , \regfile[11][7] , \regfile[11][6] ,
         \regfile[11][5] , \regfile[11][4] , \regfile[11][3] ,
         \regfile[11][2] , \regfile[11][1] , \regfile[11][0] ,
         \regfile[10][31] , \regfile[10][30] , \regfile[10][29] ,
         \regfile[10][28] , \regfile[10][27] , \regfile[10][26] ,
         \regfile[10][25] , \regfile[10][24] , \regfile[10][23] ,
         \regfile[10][22] , \regfile[10][21] , \regfile[10][20] ,
         \regfile[10][19] , \regfile[10][18] , \regfile[10][17] ,
         \regfile[10][16] , \regfile[10][15] , \regfile[10][14] ,
         \regfile[10][13] , \regfile[10][12] , \regfile[10][11] ,
         \regfile[10][10] , \regfile[10][9] , \regfile[10][8] ,
         \regfile[10][7] , \regfile[10][6] , \regfile[10][5] ,
         \regfile[10][4] , \regfile[10][3] , \regfile[10][2] ,
         \regfile[10][1] , \regfile[10][0] , \regfile[9][31] ,
         \regfile[9][30] , \regfile[9][29] , \regfile[9][28] ,
         \regfile[9][27] , \regfile[9][26] , \regfile[9][25] ,
         \regfile[9][24] , \regfile[9][23] , \regfile[9][22] ,
         \regfile[9][21] , \regfile[9][20] , \regfile[9][19] ,
         \regfile[9][18] , \regfile[9][17] , \regfile[9][16] ,
         \regfile[9][15] , \regfile[9][14] , \regfile[9][13] ,
         \regfile[9][12] , \regfile[9][11] , \regfile[9][10] , \regfile[9][9] ,
         \regfile[9][8] , \regfile[9][7] , \regfile[9][6] , \regfile[9][5] ,
         \regfile[9][4] , \regfile[9][3] , \regfile[9][2] , \regfile[9][1] ,
         \regfile[9][0] , \regfile[8][31] , \regfile[8][30] , \regfile[8][29] ,
         \regfile[8][28] , \regfile[8][27] , \regfile[8][26] ,
         \regfile[8][25] , \regfile[8][24] , \regfile[8][23] ,
         \regfile[8][22] , \regfile[8][21] , \regfile[8][20] ,
         \regfile[8][19] , \regfile[8][18] , \regfile[8][17] ,
         \regfile[8][16] , \regfile[8][15] , \regfile[8][14] ,
         \regfile[8][13] , \regfile[8][12] , \regfile[8][11] ,
         \regfile[8][10] , \regfile[8][9] , \regfile[8][8] , \regfile[8][7] ,
         \regfile[8][6] , \regfile[8][5] , \regfile[8][4] , \regfile[8][3] ,
         \regfile[8][2] , \regfile[8][1] , \regfile[8][0] , \regfile[7][31] ,
         \regfile[7][30] , \regfile[7][29] , \regfile[7][28] ,
         \regfile[7][27] , \regfile[7][26] , \regfile[7][25] ,
         \regfile[7][24] , \regfile[7][23] , \regfile[7][22] ,
         \regfile[7][21] , \regfile[7][20] , \regfile[7][19] ,
         \regfile[7][18] , \regfile[7][17] , \regfile[7][16] ,
         \regfile[7][15] , \regfile[7][14] , \regfile[7][13] ,
         \regfile[7][12] , \regfile[7][11] , \regfile[7][10] , \regfile[7][9] ,
         \regfile[7][8] , \regfile[7][7] , \regfile[7][6] , \regfile[7][5] ,
         \regfile[7][4] , \regfile[7][3] , \regfile[7][2] , \regfile[7][1] ,
         \regfile[7][0] , \regfile[6][31] , \regfile[6][30] , \regfile[6][29] ,
         \regfile[6][28] , \regfile[6][27] , \regfile[6][26] ,
         \regfile[6][25] , \regfile[6][24] , \regfile[6][23] ,
         \regfile[6][22] , \regfile[6][21] , \regfile[6][20] ,
         \regfile[6][19] , \regfile[6][18] , \regfile[6][17] ,
         \regfile[6][16] , \regfile[6][15] , \regfile[6][14] ,
         \regfile[6][13] , \regfile[6][12] , \regfile[6][11] ,
         \regfile[6][10] , \regfile[6][9] , \regfile[6][8] , \regfile[6][7] ,
         \regfile[6][6] , \regfile[6][5] , \regfile[6][4] , \regfile[6][3] ,
         \regfile[6][2] , \regfile[6][1] , \regfile[6][0] , \regfile[5][31] ,
         \regfile[5][30] , \regfile[5][29] , \regfile[5][28] ,
         \regfile[5][27] , \regfile[5][26] , \regfile[5][25] ,
         \regfile[5][24] , \regfile[5][23] , \regfile[5][22] ,
         \regfile[5][21] , \regfile[5][20] , \regfile[5][19] ,
         \regfile[5][18] , \regfile[5][17] , \regfile[5][16] ,
         \regfile[5][15] , \regfile[5][14] , \regfile[5][13] ,
         \regfile[5][12] , \regfile[5][11] , \regfile[5][10] , \regfile[5][9] ,
         \regfile[5][8] , \regfile[5][7] , \regfile[5][6] , \regfile[5][5] ,
         \regfile[5][4] , \regfile[5][3] , \regfile[5][2] , \regfile[5][1] ,
         \regfile[5][0] , \regfile[4][31] , \regfile[4][30] , \regfile[4][29] ,
         \regfile[4][28] , \regfile[4][27] , \regfile[4][26] ,
         \regfile[4][25] , \regfile[4][24] , \regfile[4][23] ,
         \regfile[4][22] , \regfile[4][21] , \regfile[4][20] ,
         \regfile[4][19] , \regfile[4][18] , \regfile[4][17] ,
         \regfile[4][16] , \regfile[4][15] , \regfile[4][14] ,
         \regfile[4][13] , \regfile[4][12] , \regfile[4][11] ,
         \regfile[4][10] , \regfile[4][9] , \regfile[4][8] , \regfile[4][7] ,
         \regfile[4][6] , \regfile[4][5] , \regfile[4][4] , \regfile[4][3] ,
         \regfile[4][2] , \regfile[4][1] , \regfile[4][0] , \regfile[3][31] ,
         \regfile[3][30] , \regfile[3][29] , \regfile[3][28] ,
         \regfile[3][27] , \regfile[3][26] , \regfile[3][25] ,
         \regfile[3][24] , \regfile[3][23] , \regfile[3][22] ,
         \regfile[3][21] , \regfile[3][20] , \regfile[3][19] ,
         \regfile[3][18] , \regfile[3][17] , \regfile[3][16] ,
         \regfile[3][15] , \regfile[3][14] , \regfile[3][13] ,
         \regfile[3][12] , \regfile[3][11] , \regfile[3][10] , \regfile[3][9] ,
         \regfile[3][8] , \regfile[3][7] , \regfile[3][6] , \regfile[3][5] ,
         \regfile[3][4] , \regfile[3][3] , \regfile[3][2] , \regfile[3][1] ,
         \regfile[3][0] , \regfile[2][31] , \regfile[2][30] , \regfile[2][29] ,
         \regfile[2][28] , \regfile[2][27] , \regfile[2][26] ,
         \regfile[2][25] , \regfile[2][24] , \regfile[2][23] ,
         \regfile[2][22] , \regfile[2][21] , \regfile[2][20] ,
         \regfile[2][19] , \regfile[2][18] , \regfile[2][17] ,
         \regfile[2][16] , \regfile[2][15] , \regfile[2][14] ,
         \regfile[2][13] , \regfile[2][12] , \regfile[2][11] ,
         \regfile[2][10] , \regfile[2][9] , \regfile[2][8] , \regfile[2][7] ,
         \regfile[2][6] , \regfile[2][5] , \regfile[2][4] , \regfile[2][3] ,
         \regfile[2][2] , \regfile[2][1] , \regfile[2][0] , \regfile[1][31] ,
         \regfile[1][30] , \regfile[1][29] , \regfile[1][28] ,
         \regfile[1][27] , \regfile[1][26] , \regfile[1][25] ,
         \regfile[1][24] , \regfile[1][23] , \regfile[1][22] ,
         \regfile[1][21] , \regfile[1][20] , \regfile[1][19] ,
         \regfile[1][18] , \regfile[1][17] , \regfile[1][16] ,
         \regfile[1][15] , \regfile[1][14] , \regfile[1][13] ,
         \regfile[1][12] , \regfile[1][11] , \regfile[1][10] , \regfile[1][9] ,
         \regfile[1][8] , \regfile[1][7] , \regfile[1][6] , \regfile[1][5] ,
         \regfile[1][4] , \regfile[1][3] , \regfile[1][2] , \regfile[1][1] ,
         \regfile[1][0] , \regfile[0][31] , \regfile[0][30] , \regfile[0][29] ,
         \regfile[0][28] , \regfile[0][27] , \regfile[0][26] ,
         \regfile[0][25] , \regfile[0][24] , \regfile[0][23] ,
         \regfile[0][22] , \regfile[0][21] , \regfile[0][20] ,
         \regfile[0][19] , \regfile[0][18] , \regfile[0][17] ,
         \regfile[0][16] , \regfile[0][15] , \regfile[0][14] ,
         \regfile[0][13] , \regfile[0][12] , \regfile[0][11] ,
         \regfile[0][10] , \regfile[0][9] , \regfile[0][8] , \regfile[0][7] ,
         \regfile[0][6] , \regfile[0][5] , \regfile[0][4] , \regfile[0][3] ,
         \regfile[0][2] , \regfile[0][1] , \regfile[0][0] , N24, N25, N26, N27,
         N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41,
         N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N324, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n314, n316, n317, n345, n346, n351, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
  wire   [31:0] IFID_A;
  wire   [31:0] IFID_B;
  wire   [3:0] IFID_dest;
  assign N15 = instr[8];
  assign N16 = instr[9];
  assign N17 = instr[10];
  assign N18 = instr[11];
  assign N19 = instr[4];
  assign N20 = instr[5];
  assign N21 = instr[6];
  assign N22 = instr[7];

  DFFX1 Carryout_reg ( .D(n1493), .CLK(clk), .Q(Carryout) );
  DFFX1 \EX_dest_reg[3]  ( .D(IFID_dest[3]), .CLK(clk), .Q(n1491) );
  DFFX1 \EX_dest_reg[2]  ( .D(IFID_dest[2]), .CLK(clk), .Q(n1489) );
  DFFX1 \EX_dest_reg[1]  ( .D(IFID_dest[1]), .CLK(clk), .Q(n1492), .QN(n1006)
         );
  DFFX1 \EX_dest_reg[0]  ( .D(IFID_dest[0]), .CLK(clk), .Q(n1490), .QN(n1007)
         );
  DFFX1 Overflow_reg ( .D(N324), .CLK(clk), .Q(Overflow) );
  DFFX1 \IFID_B_reg[31]  ( .D(n998), .CLK(clk), .Q(IFID_B[31]), .QN(n382) );
  DFFX1 \IFID_B_reg[30]  ( .D(n997), .CLK(clk), .Q(IFID_B[30]), .QN(n381) );
  DFFX1 \IFID_B_reg[29]  ( .D(n996), .CLK(clk), .Q(IFID_B[29]), .QN(n380) );
  DFFX1 \IFID_B_reg[28]  ( .D(n995), .CLK(clk), .Q(IFID_B[28]), .QN(n379) );
  DFFX1 \IFID_B_reg[27]  ( .D(n994), .CLK(clk), .Q(IFID_B[27]), .QN(n378) );
  DFFX1 \IFID_B_reg[26]  ( .D(n993), .CLK(clk), .Q(IFID_B[26]), .QN(n377) );
  DFFX1 \IFID_B_reg[25]  ( .D(n992), .CLK(clk), .Q(IFID_B[25]), .QN(n376) );
  DFFX1 \IFID_B_reg[24]  ( .D(n991), .CLK(clk), .Q(IFID_B[24]), .QN(n375) );
  DFFX1 \IFID_B_reg[23]  ( .D(n990), .CLK(clk), .Q(IFID_B[23]), .QN(n374) );
  DFFX1 \IFID_B_reg[22]  ( .D(n989), .CLK(clk), .Q(IFID_B[22]), .QN(n373) );
  DFFX1 \IFID_B_reg[21]  ( .D(n988), .CLK(clk), .Q(IFID_B[21]), .QN(n372) );
  DFFX1 \IFID_B_reg[20]  ( .D(n987), .CLK(clk), .Q(IFID_B[20]), .QN(n371) );
  DFFX1 \IFID_B_reg[19]  ( .D(n986), .CLK(clk), .Q(IFID_B[19]), .QN(n370) );
  DFFX1 \IFID_B_reg[18]  ( .D(n985), .CLK(clk), .Q(IFID_B[18]), .QN(n369) );
  DFFX1 \IFID_B_reg[17]  ( .D(n984), .CLK(clk), .Q(IFID_B[17]), .QN(n368) );
  DFFX1 \IFID_B_reg[16]  ( .D(n983), .CLK(clk), .Q(IFID_B[16]), .QN(n367) );
  DFFX1 \IFID_B_reg[15]  ( .D(n982), .CLK(clk), .Q(IFID_B[15]), .QN(n366) );
  DFFX1 \IFID_B_reg[14]  ( .D(n981), .CLK(clk), .Q(IFID_B[14]), .QN(n365) );
  DFFX1 \IFID_B_reg[13]  ( .D(n980), .CLK(clk), .Q(IFID_B[13]), .QN(n364) );
  DFFX1 \IFID_B_reg[12]  ( .D(n979), .CLK(clk), .Q(IFID_B[12]), .QN(n363) );
  DFFX1 \IFID_B_reg[11]  ( .D(n978), .CLK(clk), .Q(IFID_B[11]), .QN(n362) );
  DFFX1 \IFID_B_reg[10]  ( .D(n977), .CLK(clk), .Q(IFID_B[10]), .QN(n361) );
  DFFX1 \IFID_B_reg[9]  ( .D(n976), .CLK(clk), .Q(IFID_B[9]), .QN(n360) );
  DFFX1 \IFID_B_reg[8]  ( .D(n975), .CLK(clk), .Q(IFID_B[8]), .QN(n359) );
  DFFX1 \IFID_B_reg[7]  ( .D(n974), .CLK(clk), .Q(IFID_B[7]), .QN(n358) );
  DFFX1 \IFID_B_reg[6]  ( .D(n973), .CLK(clk), .Q(IFID_B[6]), .QN(n357) );
  DFFX1 \IFID_B_reg[5]  ( .D(n972), .CLK(clk), .Q(IFID_B[5]), .QN(n356) );
  DFFX1 \IFID_B_reg[4]  ( .D(n971), .CLK(clk), .Q(IFID_B[4]), .QN(n355) );
  DFFX1 \IFID_B_reg[3]  ( .D(n970), .CLK(clk), .Q(IFID_B[3]), .QN(n354) );
  DFFX1 \IFID_B_reg[2]  ( .D(n969), .CLK(clk), .Q(IFID_B[2]), .QN(n353) );
  DFFX1 \IFID_B_reg[1]  ( .D(n968), .CLK(clk), .Q(IFID_B[1]) );
  DFFX1 \IFID_B_reg[0]  ( .D(n967), .CLK(clk), .Q(IFID_B[0]), .QN(n351) );
  DFFX1 \IFID_ALU_ctl_reg[3]  ( .D(n966), .CLK(clk), .Q(n1488), .QN(n1003) );
  DFFX1 \IFID_ALU_ctl_reg[2]  ( .D(n965), .CLK(clk), .Q(n1487), .QN(n1001) );
  DFFX1 \IFID_ALU_ctl_reg[1]  ( .D(n964), .CLK(clk), .Q(n1486), .QN(n1005) );
  DFFX1 \IFID_ALU_ctl_reg[0]  ( .D(n963), .CLK(clk), .Q(n1485), .QN(n1002) );
  DFFX1 \IFID_A_reg[31]  ( .D(n962), .CLK(clk), .Q(IFID_A[31]), .QN(n346) );
  DFFX1 \IFID_A_reg[30]  ( .D(n961), .CLK(clk), .Q(IFID_A[30]), .QN(n345) );
  DFFX1 \IFID_A_reg[29]  ( .D(n960), .CLK(clk), .Q(IFID_A[29]) );
  DFFX1 \IFID_A_reg[28]  ( .D(n959), .CLK(clk), .Q(IFID_A[28]) );
  DFFX1 \IFID_A_reg[27]  ( .D(n958), .CLK(clk), .Q(IFID_A[27]) );
  DFFX1 \IFID_A_reg[26]  ( .D(n957), .CLK(clk), .Q(IFID_A[26]) );
  DFFX1 \IFID_A_reg[25]  ( .D(n956), .CLK(clk), .Q(IFID_A[25]) );
  DFFX1 \IFID_A_reg[24]  ( .D(n955), .CLK(clk), .Q(IFID_A[24]) );
  DFFX1 \IFID_A_reg[23]  ( .D(n954), .CLK(clk), .Q(IFID_A[23]) );
  DFFX1 \IFID_A_reg[22]  ( .D(n953), .CLK(clk), .Q(IFID_A[22]) );
  DFFX1 \IFID_A_reg[21]  ( .D(n952), .CLK(clk), .Q(IFID_A[21]) );
  DFFX1 \IFID_A_reg[20]  ( .D(n951), .CLK(clk), .Q(IFID_A[20]) );
  DFFX1 \IFID_A_reg[19]  ( .D(n950), .CLK(clk), .Q(IFID_A[19]) );
  DFFX1 \IFID_A_reg[18]  ( .D(n949), .CLK(clk), .Q(IFID_A[18]) );
  DFFX1 \IFID_A_reg[17]  ( .D(n948), .CLK(clk), .Q(IFID_A[17]) );
  DFFX1 \IFID_A_reg[16]  ( .D(n947), .CLK(clk), .Q(IFID_A[16]) );
  DFFX1 \IFID_A_reg[15]  ( .D(n946), .CLK(clk), .Q(IFID_A[15]) );
  DFFX1 \IFID_A_reg[14]  ( .D(n945), .CLK(clk), .Q(IFID_A[14]) );
  DFFX1 \IFID_A_reg[13]  ( .D(n944), .CLK(clk), .Q(IFID_A[13]) );
  DFFX1 \IFID_A_reg[12]  ( .D(n943), .CLK(clk), .Q(IFID_A[12]) );
  DFFX1 \IFID_A_reg[11]  ( .D(n942), .CLK(clk), .Q(IFID_A[11]) );
  DFFX1 \IFID_A_reg[10]  ( .D(n941), .CLK(clk), .Q(IFID_A[10]) );
  DFFX1 \IFID_A_reg[9]  ( .D(n940), .CLK(clk), .Q(IFID_A[9]) );
  DFFX1 \IFID_A_reg[8]  ( .D(n939), .CLK(clk), .Q(IFID_A[8]) );
  DFFX1 \IFID_A_reg[7]  ( .D(n938), .CLK(clk), .Q(IFID_A[7]) );
  DFFX1 \IFID_A_reg[6]  ( .D(n937), .CLK(clk), .Q(IFID_A[6]) );
  DFFX1 \IFID_A_reg[5]  ( .D(n936), .CLK(clk), .Q(IFID_A[5]) );
  DFFX1 \IFID_A_reg[4]  ( .D(n935), .CLK(clk), .Q(IFID_A[4]) );
  DFFX1 \IFID_A_reg[3]  ( .D(n934), .CLK(clk), .Q(IFID_A[3]) );
  DFFX1 \IFID_A_reg[2]  ( .D(n933), .CLK(clk), .Q(IFID_A[2]), .QN(n317) );
  DFFX1 \IFID_A_reg[1]  ( .D(n932), .CLK(clk), .Q(IFID_A[1]), .QN(n316) );
  DFFX1 \IFID_A_reg[0]  ( .D(n931), .CLK(clk), .Q(IFID_A[0]) );
  DFFX1 \IFID_dest_reg[3]  ( .D(n930), .CLK(clk), .Q(IFID_dest[3]) );
  DFFX1 \IFID_dest_reg[2]  ( .D(n929), .CLK(clk), .Q(IFID_dest[2]) );
  DFFX1 \IFID_dest_reg[1]  ( .D(n928), .CLK(clk), .Q(IFID_dest[1]) );
  DFFX1 \IFID_dest_reg[0]  ( .D(n927), .CLK(clk), .Q(IFID_dest[0]) );
  DFFX1 \AluOut_reg[31]  ( .D(n926), .CLK(clk), .Q(AluOut[31]), .QN(n314) );
  DFFARX1 \regfile_reg[0][31]  ( .D(n925), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][31] ) );
  DFFARX1 \regfile_reg[1][31]  ( .D(n924), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][31] ) );
  DFFARX1 \regfile_reg[2][31]  ( .D(n923), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][31] ) );
  DFFARX1 \regfile_reg[3][31]  ( .D(n922), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][31] ) );
  DFFARX1 \regfile_reg[4][31]  ( .D(n921), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][31] ) );
  DFFARX1 \regfile_reg[5][31]  ( .D(n920), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][31] ) );
  DFFARX1 \regfile_reg[6][31]  ( .D(n919), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][31] ) );
  DFFARX1 \regfile_reg[7][31]  ( .D(n918), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][31] ) );
  DFFARX1 \regfile_reg[8][31]  ( .D(n917), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][31] ) );
  DFFARX1 \regfile_reg[9][31]  ( .D(n916), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][31] ) );
  DFFARX1 \regfile_reg[10][31]  ( .D(n915), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][31] ) );
  DFFARX1 \regfile_reg[11][31]  ( .D(n914), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][31] ) );
  DFFARX1 \regfile_reg[12][31]  ( .D(n913), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][31] ) );
  DFFARX1 \regfile_reg[13][31]  ( .D(n912), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][31] ) );
  DFFARX1 \regfile_reg[14][31]  ( .D(n911), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][31] ) );
  DFFARX1 \regfile_reg[15][31]  ( .D(n910), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][31] ) );
  DFFX1 \AluOut_reg[30]  ( .D(n909), .CLK(clk), .Q(AluOut[30]), .QN(n309) );
  DFFARX1 \regfile_reg[0][30]  ( .D(n908), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][30] ) );
  DFFARX1 \regfile_reg[1][30]  ( .D(n907), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][30] ) );
  DFFARX1 \regfile_reg[2][30]  ( .D(n906), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][30] ) );
  DFFARX1 \regfile_reg[3][30]  ( .D(n905), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][30] ) );
  DFFARX1 \regfile_reg[4][30]  ( .D(n904), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][30] ) );
  DFFARX1 \regfile_reg[5][30]  ( .D(n903), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][30] ) );
  DFFARX1 \regfile_reg[6][30]  ( .D(n902), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][30] ) );
  DFFARX1 \regfile_reg[7][30]  ( .D(n901), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][30] ) );
  DFFARX1 \regfile_reg[8][30]  ( .D(n900), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][30] ) );
  DFFARX1 \regfile_reg[9][30]  ( .D(n899), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][30] ) );
  DFFARX1 \regfile_reg[10][30]  ( .D(n898), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][30] ) );
  DFFARX1 \regfile_reg[11][30]  ( .D(n897), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][30] ) );
  DFFARX1 \regfile_reg[12][30]  ( .D(n896), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][30] ) );
  DFFARX1 \regfile_reg[13][30]  ( .D(n895), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][30] ) );
  DFFARX1 \regfile_reg[14][30]  ( .D(n894), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][30] ) );
  DFFARX1 \regfile_reg[15][30]  ( .D(n893), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][30] ) );
  DFFX1 \AluOut_reg[29]  ( .D(n892), .CLK(clk), .Q(AluOut[29]), .QN(n308) );
  DFFARX1 \regfile_reg[0][29]  ( .D(n891), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][29] ) );
  DFFARX1 \regfile_reg[1][29]  ( .D(n890), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][29] ) );
  DFFARX1 \regfile_reg[2][29]  ( .D(n889), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][29] ) );
  DFFARX1 \regfile_reg[3][29]  ( .D(n888), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][29] ) );
  DFFARX1 \regfile_reg[4][29]  ( .D(n887), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][29] ) );
  DFFARX1 \regfile_reg[5][29]  ( .D(n886), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][29] ) );
  DFFARX1 \regfile_reg[6][29]  ( .D(n885), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][29] ) );
  DFFARX1 \regfile_reg[7][29]  ( .D(n884), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][29] ) );
  DFFARX1 \regfile_reg[8][29]  ( .D(n883), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][29] ) );
  DFFARX1 \regfile_reg[9][29]  ( .D(n882), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][29] ) );
  DFFARX1 \regfile_reg[10][29]  ( .D(n881), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][29] ) );
  DFFARX1 \regfile_reg[11][29]  ( .D(n880), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][29] ) );
  DFFARX1 \regfile_reg[12][29]  ( .D(n879), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][29] ) );
  DFFARX1 \regfile_reg[13][29]  ( .D(n878), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][29] ) );
  DFFARX1 \regfile_reg[14][29]  ( .D(n877), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][29] ) );
  DFFARX1 \regfile_reg[15][29]  ( .D(n876), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][29] ) );
  DFFX1 \AluOut_reg[28]  ( .D(n875), .CLK(clk), .Q(AluOut[28]), .QN(n307) );
  DFFARX1 \regfile_reg[0][28]  ( .D(n874), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][28] ) );
  DFFARX1 \regfile_reg[1][28]  ( .D(n873), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][28] ) );
  DFFARX1 \regfile_reg[2][28]  ( .D(n872), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][28] ) );
  DFFARX1 \regfile_reg[3][28]  ( .D(n871), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][28] ) );
  DFFARX1 \regfile_reg[4][28]  ( .D(n870), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][28] ) );
  DFFARX1 \regfile_reg[5][28]  ( .D(n869), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][28] ) );
  DFFARX1 \regfile_reg[6][28]  ( .D(n868), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][28] ) );
  DFFARX1 \regfile_reg[7][28]  ( .D(n867), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][28] ) );
  DFFARX1 \regfile_reg[8][28]  ( .D(n866), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][28] ) );
  DFFARX1 \regfile_reg[9][28]  ( .D(n865), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][28] ) );
  DFFARX1 \regfile_reg[10][28]  ( .D(n864), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][28] ) );
  DFFARX1 \regfile_reg[11][28]  ( .D(n863), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][28] ) );
  DFFARX1 \regfile_reg[12][28]  ( .D(n862), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][28] ) );
  DFFARX1 \regfile_reg[13][28]  ( .D(n861), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][28] ) );
  DFFARX1 \regfile_reg[14][28]  ( .D(n860), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][28] ) );
  DFFARX1 \regfile_reg[15][28]  ( .D(n859), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][28] ) );
  DFFX1 \AluOut_reg[27]  ( .D(n858), .CLK(clk), .Q(AluOut[27]), .QN(n306) );
  DFFARX1 \regfile_reg[0][27]  ( .D(n857), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][27] ) );
  DFFARX1 \regfile_reg[1][27]  ( .D(n856), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][27] ) );
  DFFARX1 \regfile_reg[2][27]  ( .D(n855), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][27] ) );
  DFFARX1 \regfile_reg[3][27]  ( .D(n854), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][27] ) );
  DFFARX1 \regfile_reg[4][27]  ( .D(n853), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][27] ) );
  DFFARX1 \regfile_reg[5][27]  ( .D(n852), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][27] ) );
  DFFARX1 \regfile_reg[6][27]  ( .D(n851), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][27] ) );
  DFFARX1 \regfile_reg[7][27]  ( .D(n850), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][27] ) );
  DFFARX1 \regfile_reg[8][27]  ( .D(n849), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][27] ) );
  DFFARX1 \regfile_reg[9][27]  ( .D(n848), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][27] ) );
  DFFARX1 \regfile_reg[10][27]  ( .D(n847), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][27] ) );
  DFFARX1 \regfile_reg[11][27]  ( .D(n846), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][27] ) );
  DFFARX1 \regfile_reg[12][27]  ( .D(n845), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][27] ) );
  DFFARX1 \regfile_reg[13][27]  ( .D(n844), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][27] ) );
  DFFARX1 \regfile_reg[14][27]  ( .D(n843), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][27] ) );
  DFFARX1 \regfile_reg[15][27]  ( .D(n842), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][27] ) );
  DFFX1 \AluOut_reg[26]  ( .D(n841), .CLK(clk), .Q(AluOut[26]), .QN(n305) );
  DFFARX1 \regfile_reg[0][26]  ( .D(n840), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][26] ) );
  DFFARX1 \regfile_reg[1][26]  ( .D(n839), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][26] ) );
  DFFARX1 \regfile_reg[2][26]  ( .D(n838), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][26] ) );
  DFFARX1 \regfile_reg[3][26]  ( .D(n837), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][26] ) );
  DFFARX1 \regfile_reg[4][26]  ( .D(n836), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][26] ) );
  DFFARX1 \regfile_reg[5][26]  ( .D(n835), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][26] ) );
  DFFARX1 \regfile_reg[6][26]  ( .D(n834), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][26] ) );
  DFFARX1 \regfile_reg[7][26]  ( .D(n833), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][26] ) );
  DFFARX1 \regfile_reg[8][26]  ( .D(n832), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][26] ) );
  DFFARX1 \regfile_reg[9][26]  ( .D(n831), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][26] ) );
  DFFARX1 \regfile_reg[10][26]  ( .D(n830), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][26] ) );
  DFFARX1 \regfile_reg[11][26]  ( .D(n829), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][26] ) );
  DFFARX1 \regfile_reg[12][26]  ( .D(n828), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][26] ) );
  DFFARX1 \regfile_reg[13][26]  ( .D(n827), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][26] ) );
  DFFARX1 \regfile_reg[14][26]  ( .D(n826), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][26] ) );
  DFFARX1 \regfile_reg[15][26]  ( .D(n825), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][26] ) );
  DFFX1 \AluOut_reg[25]  ( .D(n824), .CLK(clk), .Q(AluOut[25]), .QN(n304) );
  DFFARX1 \regfile_reg[0][25]  ( .D(n823), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][25] ) );
  DFFARX1 \regfile_reg[1][25]  ( .D(n822), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][25] ) );
  DFFARX1 \regfile_reg[2][25]  ( .D(n821), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][25] ) );
  DFFARX1 \regfile_reg[3][25]  ( .D(n820), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][25] ) );
  DFFARX1 \regfile_reg[4][25]  ( .D(n819), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][25] ) );
  DFFARX1 \regfile_reg[5][25]  ( .D(n818), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][25] ) );
  DFFARX1 \regfile_reg[6][25]  ( .D(n817), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][25] ) );
  DFFARX1 \regfile_reg[7][25]  ( .D(n816), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][25] ) );
  DFFARX1 \regfile_reg[8][25]  ( .D(n815), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][25] ) );
  DFFARX1 \regfile_reg[9][25]  ( .D(n814), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][25] ) );
  DFFARX1 \regfile_reg[10][25]  ( .D(n813), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][25] ) );
  DFFARX1 \regfile_reg[11][25]  ( .D(n812), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][25] ) );
  DFFARX1 \regfile_reg[12][25]  ( .D(n811), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][25] ) );
  DFFARX1 \regfile_reg[13][25]  ( .D(n810), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][25] ) );
  DFFARX1 \regfile_reg[14][25]  ( .D(n809), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][25] ) );
  DFFARX1 \regfile_reg[15][25]  ( .D(n808), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][25] ) );
  DFFX1 \AluOut_reg[24]  ( .D(n807), .CLK(clk), .Q(AluOut[24]), .QN(n303) );
  DFFARX1 \regfile_reg[0][24]  ( .D(n806), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][24] ) );
  DFFARX1 \regfile_reg[1][24]  ( .D(n805), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][24] ) );
  DFFARX1 \regfile_reg[2][24]  ( .D(n804), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][24] ) );
  DFFARX1 \regfile_reg[3][24]  ( .D(n803), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][24] ) );
  DFFARX1 \regfile_reg[4][24]  ( .D(n802), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][24] ) );
  DFFARX1 \regfile_reg[5][24]  ( .D(n801), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][24] ) );
  DFFARX1 \regfile_reg[6][24]  ( .D(n800), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][24] ) );
  DFFARX1 \regfile_reg[7][24]  ( .D(n799), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][24] ) );
  DFFARX1 \regfile_reg[8][24]  ( .D(n798), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][24] ) );
  DFFARX1 \regfile_reg[9][24]  ( .D(n797), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][24] ) );
  DFFARX1 \regfile_reg[10][24]  ( .D(n796), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][24] ) );
  DFFARX1 \regfile_reg[11][24]  ( .D(n795), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][24] ) );
  DFFARX1 \regfile_reg[12][24]  ( .D(n794), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][24] ) );
  DFFARX1 \regfile_reg[13][24]  ( .D(n793), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][24] ) );
  DFFARX1 \regfile_reg[14][24]  ( .D(n792), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][24] ) );
  DFFARX1 \regfile_reg[15][24]  ( .D(n791), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][24] ) );
  DFFX1 \AluOut_reg[23]  ( .D(n790), .CLK(clk), .Q(AluOut[23]), .QN(n302) );
  DFFARX1 \regfile_reg[0][23]  ( .D(n789), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][23] ) );
  DFFARX1 \regfile_reg[1][23]  ( .D(n788), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][23] ) );
  DFFARX1 \regfile_reg[2][23]  ( .D(n787), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][23] ) );
  DFFARX1 \regfile_reg[3][23]  ( .D(n786), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][23] ) );
  DFFARX1 \regfile_reg[4][23]  ( .D(n785), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][23] ) );
  DFFARX1 \regfile_reg[5][23]  ( .D(n784), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][23] ) );
  DFFARX1 \regfile_reg[6][23]  ( .D(n783), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][23] ) );
  DFFARX1 \regfile_reg[7][23]  ( .D(n782), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][23] ) );
  DFFARX1 \regfile_reg[8][23]  ( .D(n781), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][23] ) );
  DFFARX1 \regfile_reg[9][23]  ( .D(n780), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][23] ) );
  DFFARX1 \regfile_reg[10][23]  ( .D(n779), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][23] ) );
  DFFARX1 \regfile_reg[11][23]  ( .D(n778), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][23] ) );
  DFFARX1 \regfile_reg[12][23]  ( .D(n777), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][23] ) );
  DFFARX1 \regfile_reg[13][23]  ( .D(n776), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][23] ) );
  DFFARX1 \regfile_reg[14][23]  ( .D(n775), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][23] ) );
  DFFARX1 \regfile_reg[15][23]  ( .D(n774), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][23] ) );
  DFFX1 \AluOut_reg[22]  ( .D(n773), .CLK(clk), .Q(AluOut[22]), .QN(n301) );
  DFFARX1 \regfile_reg[0][22]  ( .D(n772), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][22] ) );
  DFFARX1 \regfile_reg[1][22]  ( .D(n771), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][22] ) );
  DFFARX1 \regfile_reg[2][22]  ( .D(n770), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][22] ) );
  DFFARX1 \regfile_reg[3][22]  ( .D(n769), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][22] ) );
  DFFARX1 \regfile_reg[4][22]  ( .D(n768), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][22] ) );
  DFFARX1 \regfile_reg[5][22]  ( .D(n767), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][22] ) );
  DFFARX1 \regfile_reg[6][22]  ( .D(n766), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][22] ) );
  DFFARX1 \regfile_reg[7][22]  ( .D(n765), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][22] ) );
  DFFARX1 \regfile_reg[8][22]  ( .D(n764), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][22] ) );
  DFFARX1 \regfile_reg[9][22]  ( .D(n763), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][22] ) );
  DFFARX1 \regfile_reg[10][22]  ( .D(n762), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][22] ) );
  DFFARX1 \regfile_reg[11][22]  ( .D(n761), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][22] ) );
  DFFARX1 \regfile_reg[12][22]  ( .D(n760), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][22] ) );
  DFFARX1 \regfile_reg[13][22]  ( .D(n759), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][22] ) );
  DFFARX1 \regfile_reg[14][22]  ( .D(n758), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][22] ) );
  DFFARX1 \regfile_reg[15][22]  ( .D(n757), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][22] ) );
  DFFX1 \AluOut_reg[21]  ( .D(n756), .CLK(clk), .Q(AluOut[21]), .QN(n300) );
  DFFARX1 \regfile_reg[0][21]  ( .D(n755), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][21] ) );
  DFFARX1 \regfile_reg[1][21]  ( .D(n754), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][21] ) );
  DFFARX1 \regfile_reg[2][21]  ( .D(n753), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][21] ) );
  DFFARX1 \regfile_reg[3][21]  ( .D(n752), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][21] ) );
  DFFARX1 \regfile_reg[4][21]  ( .D(n751), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][21] ) );
  DFFARX1 \regfile_reg[5][21]  ( .D(n750), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][21] ) );
  DFFARX1 \regfile_reg[6][21]  ( .D(n749), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][21] ) );
  DFFARX1 \regfile_reg[7][21]  ( .D(n748), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][21] ) );
  DFFARX1 \regfile_reg[8][21]  ( .D(n747), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][21] ) );
  DFFARX1 \regfile_reg[9][21]  ( .D(n746), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][21] ) );
  DFFARX1 \regfile_reg[10][21]  ( .D(n745), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][21] ) );
  DFFARX1 \regfile_reg[11][21]  ( .D(n744), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][21] ) );
  DFFARX1 \regfile_reg[12][21]  ( .D(n743), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][21] ) );
  DFFARX1 \regfile_reg[13][21]  ( .D(n742), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][21] ) );
  DFFARX1 \regfile_reg[14][21]  ( .D(n741), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][21] ) );
  DFFARX1 \regfile_reg[15][21]  ( .D(n740), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][21] ) );
  DFFX1 \AluOut_reg[20]  ( .D(n739), .CLK(clk), .Q(AluOut[20]), .QN(n299) );
  DFFARX1 \regfile_reg[0][20]  ( .D(n738), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][20] ) );
  DFFARX1 \regfile_reg[1][20]  ( .D(n737), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][20] ) );
  DFFARX1 \regfile_reg[2][20]  ( .D(n736), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][20] ) );
  DFFARX1 \regfile_reg[3][20]  ( .D(n735), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][20] ) );
  DFFARX1 \regfile_reg[4][20]  ( .D(n734), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][20] ) );
  DFFARX1 \regfile_reg[5][20]  ( .D(n733), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][20] ) );
  DFFARX1 \regfile_reg[6][20]  ( .D(n732), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][20] ) );
  DFFARX1 \regfile_reg[7][20]  ( .D(n731), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][20] ) );
  DFFARX1 \regfile_reg[8][20]  ( .D(n730), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][20] ) );
  DFFARX1 \regfile_reg[9][20]  ( .D(n729), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][20] ) );
  DFFARX1 \regfile_reg[10][20]  ( .D(n728), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][20] ) );
  DFFARX1 \regfile_reg[11][20]  ( .D(n727), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][20] ) );
  DFFARX1 \regfile_reg[12][20]  ( .D(n726), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][20] ) );
  DFFARX1 \regfile_reg[13][20]  ( .D(n725), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][20] ) );
  DFFARX1 \regfile_reg[14][20]  ( .D(n724), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][20] ) );
  DFFARX1 \regfile_reg[15][20]  ( .D(n723), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][20] ) );
  DFFX1 \AluOut_reg[19]  ( .D(n722), .CLK(clk), .Q(AluOut[19]), .QN(n298) );
  DFFARX1 \regfile_reg[0][19]  ( .D(n721), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][19] ) );
  DFFARX1 \regfile_reg[1][19]  ( .D(n720), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][19] ) );
  DFFARX1 \regfile_reg[2][19]  ( .D(n719), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][19] ) );
  DFFARX1 \regfile_reg[3][19]  ( .D(n718), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][19] ) );
  DFFARX1 \regfile_reg[4][19]  ( .D(n717), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][19] ) );
  DFFARX1 \regfile_reg[5][19]  ( .D(n716), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][19] ) );
  DFFARX1 \regfile_reg[6][19]  ( .D(n715), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][19] ) );
  DFFARX1 \regfile_reg[7][19]  ( .D(n714), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][19] ) );
  DFFARX1 \regfile_reg[8][19]  ( .D(n713), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][19] ) );
  DFFARX1 \regfile_reg[9][19]  ( .D(n712), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][19] ) );
  DFFARX1 \regfile_reg[10][19]  ( .D(n711), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][19] ) );
  DFFARX1 \regfile_reg[11][19]  ( .D(n710), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][19] ) );
  DFFARX1 \regfile_reg[12][19]  ( .D(n709), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][19] ) );
  DFFARX1 \regfile_reg[13][19]  ( .D(n708), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][19] ) );
  DFFARX1 \regfile_reg[14][19]  ( .D(n707), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][19] ) );
  DFFARX1 \regfile_reg[15][19]  ( .D(n706), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][19] ) );
  DFFX1 \AluOut_reg[18]  ( .D(n705), .CLK(clk), .Q(AluOut[18]), .QN(n297) );
  DFFARX1 \regfile_reg[0][18]  ( .D(n704), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][18] ) );
  DFFARX1 \regfile_reg[1][18]  ( .D(n703), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][18] ) );
  DFFARX1 \regfile_reg[2][18]  ( .D(n702), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][18] ) );
  DFFARX1 \regfile_reg[3][18]  ( .D(n701), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][18] ) );
  DFFARX1 \regfile_reg[4][18]  ( .D(n700), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][18] ) );
  DFFARX1 \regfile_reg[5][18]  ( .D(n699), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][18] ) );
  DFFARX1 \regfile_reg[6][18]  ( .D(n698), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][18] ) );
  DFFARX1 \regfile_reg[7][18]  ( .D(n697), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][18] ) );
  DFFARX1 \regfile_reg[8][18]  ( .D(n696), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][18] ) );
  DFFARX1 \regfile_reg[9][18]  ( .D(n695), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][18] ) );
  DFFARX1 \regfile_reg[10][18]  ( .D(n694), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][18] ) );
  DFFARX1 \regfile_reg[11][18]  ( .D(n693), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][18] ) );
  DFFARX1 \regfile_reg[12][18]  ( .D(n692), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][18] ) );
  DFFARX1 \regfile_reg[13][18]  ( .D(n691), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][18] ) );
  DFFARX1 \regfile_reg[14][18]  ( .D(n690), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][18] ) );
  DFFARX1 \regfile_reg[15][18]  ( .D(n689), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][18] ) );
  DFFX1 \AluOut_reg[17]  ( .D(n688), .CLK(clk), .Q(AluOut[17]), .QN(n296) );
  DFFARX1 \regfile_reg[0][17]  ( .D(n687), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][17] ) );
  DFFARX1 \regfile_reg[1][17]  ( .D(n686), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][17] ) );
  DFFARX1 \regfile_reg[2][17]  ( .D(n685), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][17] ) );
  DFFARX1 \regfile_reg[3][17]  ( .D(n684), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][17] ) );
  DFFARX1 \regfile_reg[4][17]  ( .D(n683), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][17] ) );
  DFFARX1 \regfile_reg[5][17]  ( .D(n682), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][17] ) );
  DFFARX1 \regfile_reg[6][17]  ( .D(n681), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][17] ) );
  DFFARX1 \regfile_reg[7][17]  ( .D(n680), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][17] ) );
  DFFARX1 \regfile_reg[8][17]  ( .D(n679), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][17] ) );
  DFFARX1 \regfile_reg[9][17]  ( .D(n678), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][17] ) );
  DFFARX1 \regfile_reg[10][17]  ( .D(n677), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][17] ) );
  DFFARX1 \regfile_reg[11][17]  ( .D(n676), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][17] ) );
  DFFARX1 \regfile_reg[12][17]  ( .D(n675), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][17] ) );
  DFFARX1 \regfile_reg[13][17]  ( .D(n674), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][17] ) );
  DFFARX1 \regfile_reg[14][17]  ( .D(n673), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][17] ) );
  DFFARX1 \regfile_reg[15][17]  ( .D(n672), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][17] ) );
  DFFX1 \AluOut_reg[16]  ( .D(n671), .CLK(clk), .Q(AluOut[16]), .QN(n295) );
  DFFARX1 \regfile_reg[0][16]  ( .D(n670), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][16] ) );
  DFFARX1 \regfile_reg[1][16]  ( .D(n669), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][16] ) );
  DFFARX1 \regfile_reg[2][16]  ( .D(n668), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][16] ) );
  DFFARX1 \regfile_reg[3][16]  ( .D(n667), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][16] ) );
  DFFARX1 \regfile_reg[4][16]  ( .D(n666), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][16] ) );
  DFFARX1 \regfile_reg[5][16]  ( .D(n665), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][16] ) );
  DFFARX1 \regfile_reg[6][16]  ( .D(n664), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][16] ) );
  DFFARX1 \regfile_reg[7][16]  ( .D(n663), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][16] ) );
  DFFARX1 \regfile_reg[8][16]  ( .D(n662), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][16] ) );
  DFFARX1 \regfile_reg[9][16]  ( .D(n661), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][16] ) );
  DFFARX1 \regfile_reg[10][16]  ( .D(n660), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][16] ) );
  DFFARX1 \regfile_reg[11][16]  ( .D(n659), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][16] ) );
  DFFARX1 \regfile_reg[12][16]  ( .D(n658), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][16] ) );
  DFFARX1 \regfile_reg[13][16]  ( .D(n657), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][16] ) );
  DFFARX1 \regfile_reg[14][16]  ( .D(n656), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][16] ) );
  DFFARX1 \regfile_reg[15][16]  ( .D(n655), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][16] ) );
  DFFX1 \AluOut_reg[15]  ( .D(n654), .CLK(clk), .Q(AluOut[15]), .QN(n294) );
  DFFARX1 \regfile_reg[0][15]  ( .D(n653), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][15] ) );
  DFFARX1 \regfile_reg[1][15]  ( .D(n652), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][15] ) );
  DFFARX1 \regfile_reg[2][15]  ( .D(n651), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][15] ) );
  DFFARX1 \regfile_reg[3][15]  ( .D(n650), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][15] ) );
  DFFARX1 \regfile_reg[4][15]  ( .D(n649), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][15] ) );
  DFFARX1 \regfile_reg[5][15]  ( .D(n648), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][15] ) );
  DFFARX1 \regfile_reg[6][15]  ( .D(n647), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][15] ) );
  DFFARX1 \regfile_reg[7][15]  ( .D(n646), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][15] ) );
  DFFARX1 \regfile_reg[8][15]  ( .D(n645), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][15] ) );
  DFFARX1 \regfile_reg[9][15]  ( .D(n644), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][15] ) );
  DFFARX1 \regfile_reg[10][15]  ( .D(n643), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][15] ) );
  DFFARX1 \regfile_reg[11][15]  ( .D(n642), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][15] ) );
  DFFARX1 \regfile_reg[12][15]  ( .D(n641), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][15] ) );
  DFFARX1 \regfile_reg[13][15]  ( .D(n640), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][15] ) );
  DFFARX1 \regfile_reg[14][15]  ( .D(n639), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][15] ) );
  DFFARX1 \regfile_reg[15][15]  ( .D(n638), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][15] ) );
  DFFX1 \AluOut_reg[14]  ( .D(n637), .CLK(clk), .Q(AluOut[14]), .QN(n293) );
  DFFARX1 \regfile_reg[0][14]  ( .D(n636), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][14] ) );
  DFFARX1 \regfile_reg[1][14]  ( .D(n635), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][14] ) );
  DFFARX1 \regfile_reg[2][14]  ( .D(n634), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][14] ) );
  DFFARX1 \regfile_reg[3][14]  ( .D(n633), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][14] ) );
  DFFARX1 \regfile_reg[4][14]  ( .D(n632), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][14] ) );
  DFFARX1 \regfile_reg[5][14]  ( .D(n631), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][14] ) );
  DFFARX1 \regfile_reg[6][14]  ( .D(n630), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][14] ) );
  DFFARX1 \regfile_reg[7][14]  ( .D(n629), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][14] ) );
  DFFARX1 \regfile_reg[8][14]  ( .D(n628), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][14] ) );
  DFFARX1 \regfile_reg[9][14]  ( .D(n627), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][14] ) );
  DFFARX1 \regfile_reg[10][14]  ( .D(n626), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][14] ) );
  DFFARX1 \regfile_reg[11][14]  ( .D(n625), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][14] ) );
  DFFARX1 \regfile_reg[12][14]  ( .D(n624), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][14] ) );
  DFFARX1 \regfile_reg[13][14]  ( .D(n623), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][14] ) );
  DFFARX1 \regfile_reg[14][14]  ( .D(n622), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][14] ) );
  DFFARX1 \regfile_reg[15][14]  ( .D(n621), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][14] ) );
  DFFX1 \AluOut_reg[13]  ( .D(n620), .CLK(clk), .Q(AluOut[13]), .QN(n292) );
  DFFARX1 \regfile_reg[0][13]  ( .D(n619), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][13] ) );
  DFFARX1 \regfile_reg[1][13]  ( .D(n618), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][13] ) );
  DFFARX1 \regfile_reg[2][13]  ( .D(n617), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][13] ) );
  DFFARX1 \regfile_reg[3][13]  ( .D(n616), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][13] ) );
  DFFARX1 \regfile_reg[4][13]  ( .D(n615), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][13] ) );
  DFFARX1 \regfile_reg[5][13]  ( .D(n614), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][13] ) );
  DFFARX1 \regfile_reg[6][13]  ( .D(n613), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][13] ) );
  DFFARX1 \regfile_reg[7][13]  ( .D(n612), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][13] ) );
  DFFARX1 \regfile_reg[8][13]  ( .D(n611), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][13] ) );
  DFFARX1 \regfile_reg[9][13]  ( .D(n610), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][13] ) );
  DFFARX1 \regfile_reg[10][13]  ( .D(n609), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][13] ) );
  DFFARX1 \regfile_reg[11][13]  ( .D(n608), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][13] ) );
  DFFARX1 \regfile_reg[12][13]  ( .D(n607), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][13] ) );
  DFFARX1 \regfile_reg[13][13]  ( .D(n606), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][13] ) );
  DFFARX1 \regfile_reg[14][13]  ( .D(n605), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][13] ) );
  DFFARX1 \regfile_reg[15][13]  ( .D(n604), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][13] ) );
  DFFX1 \AluOut_reg[12]  ( .D(n603), .CLK(clk), .Q(AluOut[12]), .QN(n291) );
  DFFARX1 \regfile_reg[0][12]  ( .D(n602), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][12] ) );
  DFFARX1 \regfile_reg[1][12]  ( .D(n601), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][12] ) );
  DFFARX1 \regfile_reg[2][12]  ( .D(n600), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][12] ) );
  DFFARX1 \regfile_reg[3][12]  ( .D(n599), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][12] ) );
  DFFARX1 \regfile_reg[4][12]  ( .D(n598), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][12] ) );
  DFFARX1 \regfile_reg[5][12]  ( .D(n597), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][12] ) );
  DFFARX1 \regfile_reg[6][12]  ( .D(n596), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][12] ) );
  DFFARX1 \regfile_reg[7][12]  ( .D(n595), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][12] ) );
  DFFARX1 \regfile_reg[8][12]  ( .D(n594), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][12] ) );
  DFFARX1 \regfile_reg[9][12]  ( .D(n593), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][12] ) );
  DFFARX1 \regfile_reg[10][12]  ( .D(n592), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][12] ) );
  DFFARX1 \regfile_reg[11][12]  ( .D(n591), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][12] ) );
  DFFARX1 \regfile_reg[12][12]  ( .D(n590), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][12] ) );
  DFFARX1 \regfile_reg[13][12]  ( .D(n589), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][12] ) );
  DFFARX1 \regfile_reg[14][12]  ( .D(n588), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][12] ) );
  DFFARX1 \regfile_reg[15][12]  ( .D(n587), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][12] ) );
  DFFX1 \AluOut_reg[11]  ( .D(n586), .CLK(clk), .Q(AluOut[11]), .QN(n290) );
  DFFARX1 \regfile_reg[0][11]  ( .D(n585), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][11] ) );
  DFFARX1 \regfile_reg[1][11]  ( .D(n584), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][11] ) );
  DFFARX1 \regfile_reg[2][11]  ( .D(n583), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][11] ) );
  DFFARX1 \regfile_reg[3][11]  ( .D(n582), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][11] ) );
  DFFARX1 \regfile_reg[4][11]  ( .D(n581), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][11] ) );
  DFFARX1 \regfile_reg[5][11]  ( .D(n580), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][11] ) );
  DFFARX1 \regfile_reg[6][11]  ( .D(n579), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][11] ) );
  DFFARX1 \regfile_reg[7][11]  ( .D(n578), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][11] ) );
  DFFARX1 \regfile_reg[8][11]  ( .D(n577), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][11] ) );
  DFFARX1 \regfile_reg[9][11]  ( .D(n576), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][11] ) );
  DFFARX1 \regfile_reg[10][11]  ( .D(n575), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][11] ) );
  DFFARX1 \regfile_reg[11][11]  ( .D(n574), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][11] ) );
  DFFARX1 \regfile_reg[12][11]  ( .D(n573), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][11] ) );
  DFFARX1 \regfile_reg[13][11]  ( .D(n572), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][11] ) );
  DFFARX1 \regfile_reg[14][11]  ( .D(n571), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][11] ) );
  DFFARX1 \regfile_reg[15][11]  ( .D(n570), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][11] ) );
  DFFX1 \AluOut_reg[10]  ( .D(n569), .CLK(clk), .Q(AluOut[10]), .QN(n289) );
  DFFARX1 \regfile_reg[0][10]  ( .D(n568), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][10] ) );
  DFFARX1 \regfile_reg[1][10]  ( .D(n567), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][10] ) );
  DFFARX1 \regfile_reg[2][10]  ( .D(n566), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][10] ) );
  DFFARX1 \regfile_reg[3][10]  ( .D(n565), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][10] ) );
  DFFARX1 \regfile_reg[4][10]  ( .D(n564), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][10] ) );
  DFFARX1 \regfile_reg[5][10]  ( .D(n563), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][10] ) );
  DFFARX1 \regfile_reg[6][10]  ( .D(n562), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][10] ) );
  DFFARX1 \regfile_reg[7][10]  ( .D(n561), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][10] ) );
  DFFARX1 \regfile_reg[8][10]  ( .D(n560), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][10] ) );
  DFFARX1 \regfile_reg[9][10]  ( .D(n559), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][10] ) );
  DFFARX1 \regfile_reg[10][10]  ( .D(n558), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][10] ) );
  DFFARX1 \regfile_reg[11][10]  ( .D(n557), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][10] ) );
  DFFARX1 \regfile_reg[12][10]  ( .D(n556), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][10] ) );
  DFFARX1 \regfile_reg[13][10]  ( .D(n555), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][10] ) );
  DFFARX1 \regfile_reg[14][10]  ( .D(n554), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][10] ) );
  DFFARX1 \regfile_reg[15][10]  ( .D(n553), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][10] ) );
  DFFX1 \AluOut_reg[9]  ( .D(n552), .CLK(clk), .Q(AluOut[9]), .QN(n288) );
  DFFARX1 \regfile_reg[0][9]  ( .D(n551), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][9] ) );
  DFFARX1 \regfile_reg[1][9]  ( .D(n550), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][9] ) );
  DFFARX1 \regfile_reg[2][9]  ( .D(n549), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][9] ) );
  DFFARX1 \regfile_reg[3][9]  ( .D(n548), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][9] ) );
  DFFARX1 \regfile_reg[4][9]  ( .D(n547), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][9] ) );
  DFFARX1 \regfile_reg[5][9]  ( .D(n546), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][9] ) );
  DFFARX1 \regfile_reg[6][9]  ( .D(n545), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][9] ) );
  DFFARX1 \regfile_reg[7][9]  ( .D(n544), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][9] ) );
  DFFARX1 \regfile_reg[8][9]  ( .D(n543), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][9] ) );
  DFFARX1 \regfile_reg[9][9]  ( .D(n542), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][9] ) );
  DFFARX1 \regfile_reg[10][9]  ( .D(n541), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][9] ) );
  DFFARX1 \regfile_reg[11][9]  ( .D(n540), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][9] ) );
  DFFARX1 \regfile_reg[12][9]  ( .D(n539), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][9] ) );
  DFFARX1 \regfile_reg[13][9]  ( .D(n538), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][9] ) );
  DFFARX1 \regfile_reg[14][9]  ( .D(n537), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][9] ) );
  DFFARX1 \regfile_reg[15][9]  ( .D(n536), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][9] ) );
  DFFX1 \AluOut_reg[8]  ( .D(n535), .CLK(clk), .Q(AluOut[8]), .QN(n287) );
  DFFARX1 \regfile_reg[0][8]  ( .D(n534), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][8] ) );
  DFFARX1 \regfile_reg[1][8]  ( .D(n533), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][8] ) );
  DFFARX1 \regfile_reg[2][8]  ( .D(n532), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][8] ) );
  DFFARX1 \regfile_reg[3][8]  ( .D(n531), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][8] ) );
  DFFARX1 \regfile_reg[4][8]  ( .D(n530), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][8] ) );
  DFFARX1 \regfile_reg[5][8]  ( .D(n529), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][8] ) );
  DFFARX1 \regfile_reg[6][8]  ( .D(n528), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][8] ) );
  DFFARX1 \regfile_reg[7][8]  ( .D(n527), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][8] ) );
  DFFARX1 \regfile_reg[8][8]  ( .D(n526), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][8] ) );
  DFFARX1 \regfile_reg[9][8]  ( .D(n525), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][8] ) );
  DFFARX1 \regfile_reg[10][8]  ( .D(n524), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][8] ) );
  DFFARX1 \regfile_reg[11][8]  ( .D(n523), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][8] ) );
  DFFARX1 \regfile_reg[12][8]  ( .D(n522), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][8] ) );
  DFFARX1 \regfile_reg[13][8]  ( .D(n521), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][8] ) );
  DFFARX1 \regfile_reg[14][8]  ( .D(n520), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][8] ) );
  DFFARX1 \regfile_reg[15][8]  ( .D(n519), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][8] ) );
  DFFX1 \AluOut_reg[7]  ( .D(n518), .CLK(clk), .Q(AluOut[7]), .QN(n286) );
  DFFARX1 \regfile_reg[0][7]  ( .D(n517), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][7] ) );
  DFFARX1 \regfile_reg[1][7]  ( .D(n516), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][7] ) );
  DFFARX1 \regfile_reg[2][7]  ( .D(n515), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][7] ) );
  DFFARX1 \regfile_reg[3][7]  ( .D(n514), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][7] ) );
  DFFARX1 \regfile_reg[4][7]  ( .D(n513), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][7] ) );
  DFFARX1 \regfile_reg[5][7]  ( .D(n512), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][7] ) );
  DFFARX1 \regfile_reg[6][7]  ( .D(n511), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][7] ) );
  DFFARX1 \regfile_reg[7][7]  ( .D(n510), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][7] ) );
  DFFARX1 \regfile_reg[8][7]  ( .D(n509), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][7] ) );
  DFFARX1 \regfile_reg[9][7]  ( .D(n508), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][7] ) );
  DFFARX1 \regfile_reg[10][7]  ( .D(n507), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][7] ) );
  DFFARX1 \regfile_reg[11][7]  ( .D(n506), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][7] ) );
  DFFARX1 \regfile_reg[12][7]  ( .D(n505), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][7] ) );
  DFFARX1 \regfile_reg[13][7]  ( .D(n504), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][7] ) );
  DFFARX1 \regfile_reg[14][7]  ( .D(n503), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][7] ) );
  DFFARX1 \regfile_reg[15][7]  ( .D(n502), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][7] ) );
  DFFX1 \AluOut_reg[6]  ( .D(n501), .CLK(clk), .Q(AluOut[6]), .QN(n285) );
  DFFARX1 \regfile_reg[0][6]  ( .D(n500), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][6] ) );
  DFFARX1 \regfile_reg[1][6]  ( .D(n499), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][6] ) );
  DFFARX1 \regfile_reg[2][6]  ( .D(n498), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][6] ) );
  DFFARX1 \regfile_reg[3][6]  ( .D(n497), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][6] ) );
  DFFARX1 \regfile_reg[4][6]  ( .D(n496), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][6] ) );
  DFFARX1 \regfile_reg[5][6]  ( .D(n495), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][6] ) );
  DFFARX1 \regfile_reg[6][6]  ( .D(n494), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][6] ) );
  DFFARX1 \regfile_reg[7][6]  ( .D(n493), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][6] ) );
  DFFARX1 \regfile_reg[8][6]  ( .D(n492), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][6] ) );
  DFFARX1 \regfile_reg[9][6]  ( .D(n491), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][6] ) );
  DFFARX1 \regfile_reg[10][6]  ( .D(n490), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][6] ) );
  DFFARX1 \regfile_reg[11][6]  ( .D(n489), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][6] ) );
  DFFARX1 \regfile_reg[12][6]  ( .D(n488), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][6] ) );
  DFFARX1 \regfile_reg[13][6]  ( .D(n487), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][6] ) );
  DFFARX1 \regfile_reg[14][6]  ( .D(n486), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][6] ) );
  DFFARX1 \regfile_reg[15][6]  ( .D(n485), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][6] ) );
  DFFX1 \AluOut_reg[5]  ( .D(n484), .CLK(clk), .Q(AluOut[5]), .QN(n284) );
  DFFARX1 \regfile_reg[0][5]  ( .D(n483), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][5] ) );
  DFFARX1 \regfile_reg[1][5]  ( .D(n482), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][5] ) );
  DFFARX1 \regfile_reg[2][5]  ( .D(n481), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][5] ) );
  DFFARX1 \regfile_reg[3][5]  ( .D(n480), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][5] ) );
  DFFARX1 \regfile_reg[4][5]  ( .D(n479), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][5] ) );
  DFFARX1 \regfile_reg[5][5]  ( .D(n478), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][5] ) );
  DFFARX1 \regfile_reg[6][5]  ( .D(n477), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][5] ) );
  DFFARX1 \regfile_reg[7][5]  ( .D(n476), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][5] ) );
  DFFARX1 \regfile_reg[8][5]  ( .D(n475), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][5] ) );
  DFFARX1 \regfile_reg[9][5]  ( .D(n474), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][5] ) );
  DFFARX1 \regfile_reg[10][5]  ( .D(n473), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][5] ) );
  DFFARX1 \regfile_reg[11][5]  ( .D(n472), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][5] ) );
  DFFARX1 \regfile_reg[12][5]  ( .D(n471), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][5] ) );
  DFFARX1 \regfile_reg[13][5]  ( .D(n470), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][5] ) );
  DFFARX1 \regfile_reg[14][5]  ( .D(n469), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][5] ) );
  DFFARX1 \regfile_reg[15][5]  ( .D(n468), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][5] ) );
  DFFX1 \AluOut_reg[4]  ( .D(n467), .CLK(clk), .Q(AluOut[4]), .QN(n283) );
  DFFARX1 \regfile_reg[0][4]  ( .D(n466), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][4] ) );
  DFFARX1 \regfile_reg[1][4]  ( .D(n465), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][4] ) );
  DFFARX1 \regfile_reg[2][4]  ( .D(n464), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][4] ) );
  DFFARX1 \regfile_reg[3][4]  ( .D(n463), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][4] ) );
  DFFARX1 \regfile_reg[4][4]  ( .D(n462), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][4] ) );
  DFFARX1 \regfile_reg[5][4]  ( .D(n461), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][4] ) );
  DFFARX1 \regfile_reg[6][4]  ( .D(n460), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][4] ) );
  DFFARX1 \regfile_reg[7][4]  ( .D(n459), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][4] ) );
  DFFARX1 \regfile_reg[8][4]  ( .D(n458), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][4] ) );
  DFFARX1 \regfile_reg[9][4]  ( .D(n457), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][4] ) );
  DFFARX1 \regfile_reg[10][4]  ( .D(n456), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][4] ) );
  DFFARX1 \regfile_reg[11][4]  ( .D(n455), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][4] ) );
  DFFARX1 \regfile_reg[12][4]  ( .D(n454), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][4] ) );
  DFFARX1 \regfile_reg[13][4]  ( .D(n453), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][4] ) );
  DFFARX1 \regfile_reg[14][4]  ( .D(n452), .CLK(clk), .RSTB(rst), .Q(
        \regfile[14][4] ) );
  DFFASX1 \regfile_reg[15][4]  ( .D(n451), .CLK(clk), .SETB(rst), .Q(
        \regfile[15][4] ) );
  DFFX1 \AluOut_reg[3]  ( .D(n450), .CLK(clk), .Q(AluOut[3]), .QN(n282) );
  DFFARX1 \regfile_reg[0][3]  ( .D(n449), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][3] ) );
  DFFARX1 \regfile_reg[1][3]  ( .D(n448), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][3] ) );
  DFFARX1 \regfile_reg[2][3]  ( .D(n447), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][3] ) );
  DFFARX1 \regfile_reg[3][3]  ( .D(n446), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][3] ) );
  DFFARX1 \regfile_reg[4][3]  ( .D(n445), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][3] ) );
  DFFARX1 \regfile_reg[5][3]  ( .D(n444), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][3] ) );
  DFFARX1 \regfile_reg[6][3]  ( .D(n443), .CLK(clk), .RSTB(rst), .Q(
        \regfile[6][3] ) );
  DFFASX1 \regfile_reg[7][3]  ( .D(n442), .CLK(clk), .SETB(rst), .Q(
        \regfile[7][3] ) );
  DFFASX1 \regfile_reg[8][3]  ( .D(n441), .CLK(clk), .SETB(rst), .Q(
        \regfile[8][3] ) );
  DFFASX1 \regfile_reg[9][3]  ( .D(n440), .CLK(clk), .SETB(rst), .Q(
        \regfile[9][3] ) );
  DFFASX1 \regfile_reg[10][3]  ( .D(n439), .CLK(clk), .SETB(rst), .Q(
        \regfile[10][3] ) );
  DFFASX1 \regfile_reg[11][3]  ( .D(n438), .CLK(clk), .SETB(rst), .Q(
        \regfile[11][3] ) );
  DFFASX1 \regfile_reg[12][3]  ( .D(n437), .CLK(clk), .SETB(rst), .Q(
        \regfile[12][3] ) );
  DFFASX1 \regfile_reg[13][3]  ( .D(n436), .CLK(clk), .SETB(rst), .Q(
        \regfile[13][3] ) );
  DFFASX1 \regfile_reg[14][3]  ( .D(n435), .CLK(clk), .SETB(rst), .Q(
        \regfile[14][3] ) );
  DFFARX1 \regfile_reg[15][3]  ( .D(n434), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][3] ) );
  DFFX1 \AluOut_reg[2]  ( .D(n433), .CLK(clk), .Q(AluOut[2]), .QN(n281) );
  DFFARX1 \regfile_reg[0][2]  ( .D(n432), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][2] ) );
  DFFARX1 \regfile_reg[1][2]  ( .D(n431), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][2] ) );
  DFFARX1 \regfile_reg[2][2]  ( .D(n430), .CLK(clk), .RSTB(rst), .Q(
        \regfile[2][2] ) );
  DFFASX1 \regfile_reg[3][2]  ( .D(n429), .CLK(clk), .SETB(rst), .Q(
        \regfile[3][2] ) );
  DFFASX1 \regfile_reg[4][2]  ( .D(n428), .CLK(clk), .SETB(rst), .Q(
        \regfile[4][2] ) );
  DFFASX1 \regfile_reg[5][2]  ( .D(n427), .CLK(clk), .SETB(rst), .Q(
        \regfile[5][2] ) );
  DFFASX1 \regfile_reg[6][2]  ( .D(n426), .CLK(clk), .SETB(rst), .Q(
        \regfile[6][2] ) );
  DFFARX1 \regfile_reg[7][2]  ( .D(n425), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][2] ) );
  DFFARX1 \regfile_reg[8][2]  ( .D(n424), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][2] ) );
  DFFARX1 \regfile_reg[9][2]  ( .D(n423), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][2] ) );
  DFFARX1 \regfile_reg[10][2]  ( .D(n422), .CLK(clk), .RSTB(rst), .Q(
        \regfile[10][2] ) );
  DFFASX1 \regfile_reg[11][2]  ( .D(n421), .CLK(clk), .SETB(rst), .Q(
        \regfile[11][2] ) );
  DFFASX1 \regfile_reg[12][2]  ( .D(n420), .CLK(clk), .SETB(rst), .Q(
        \regfile[12][2] ) );
  DFFASX1 \regfile_reg[13][2]  ( .D(n419), .CLK(clk), .SETB(rst), .Q(
        \regfile[13][2] ) );
  DFFASX1 \regfile_reg[14][2]  ( .D(n418), .CLK(clk), .SETB(rst), .Q(
        \regfile[14][2] ) );
  DFFARX1 \regfile_reg[15][2]  ( .D(n417), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][2] ) );
  DFFX1 \AluOut_reg[1]  ( .D(n416), .CLK(clk), .Q(AluOut[1]), .QN(n280) );
  DFFARX1 \regfile_reg[0][1]  ( .D(n415), .CLK(clk), .RSTB(rst), .Q(
        \regfile[0][1] ) );
  DFFASX1 \regfile_reg[1][1]  ( .D(n414), .CLK(clk), .SETB(rst), .Q(
        \regfile[1][1] ) );
  DFFASX1 \regfile_reg[2][1]  ( .D(n413), .CLK(clk), .SETB(rst), .Q(
        \regfile[2][1] ) );
  DFFARX1 \regfile_reg[3][1]  ( .D(n412), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][1] ) );
  DFFARX1 \regfile_reg[4][1]  ( .D(n411), .CLK(clk), .RSTB(rst), .Q(
        \regfile[4][1] ) );
  DFFASX1 \regfile_reg[5][1]  ( .D(n410), .CLK(clk), .SETB(rst), .Q(
        \regfile[5][1] ) );
  DFFASX1 \regfile_reg[6][1]  ( .D(n409), .CLK(clk), .SETB(rst), .Q(
        \regfile[6][1] ) );
  DFFARX1 \regfile_reg[7][1]  ( .D(n408), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][1] ) );
  DFFARX1 \regfile_reg[8][1]  ( .D(n407), .CLK(clk), .RSTB(rst), .Q(
        \regfile[8][1] ) );
  DFFASX1 \regfile_reg[9][1]  ( .D(n406), .CLK(clk), .SETB(rst), .Q(
        \regfile[9][1] ) );
  DFFASX1 \regfile_reg[10][1]  ( .D(n405), .CLK(clk), .SETB(rst), .Q(
        \regfile[10][1] ) );
  DFFARX1 \regfile_reg[11][1]  ( .D(n404), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][1] ) );
  DFFARX1 \regfile_reg[12][1]  ( .D(n403), .CLK(clk), .RSTB(rst), .Q(
        \regfile[12][1] ) );
  DFFASX1 \regfile_reg[13][1]  ( .D(n402), .CLK(clk), .SETB(rst), .Q(
        \regfile[13][1] ) );
  DFFASX1 \regfile_reg[14][1]  ( .D(n401), .CLK(clk), .SETB(rst), .Q(
        \regfile[14][1] ) );
  DFFARX1 \regfile_reg[15][1]  ( .D(n400), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][1] ) );
  DFFX1 \AluOut_reg[0]  ( .D(n399), .CLK(clk), .Q(AluOut[0]), .QN(n279) );
  DFFASX1 \regfile_reg[0][0]  ( .D(n398), .CLK(clk), .SETB(rst), .Q(
        \regfile[0][0] ) );
  DFFARX1 \regfile_reg[1][0]  ( .D(n397), .CLK(clk), .RSTB(rst), .Q(
        \regfile[1][0] ) );
  DFFASX1 \regfile_reg[2][0]  ( .D(n396), .CLK(clk), .SETB(rst), .Q(
        \regfile[2][0] ) );
  DFFARX1 \regfile_reg[3][0]  ( .D(n395), .CLK(clk), .RSTB(rst), .Q(
        \regfile[3][0] ) );
  DFFASX1 \regfile_reg[4][0]  ( .D(n394), .CLK(clk), .SETB(rst), .Q(
        \regfile[4][0] ) );
  DFFARX1 \regfile_reg[5][0]  ( .D(n393), .CLK(clk), .RSTB(rst), .Q(
        \regfile[5][0] ) );
  DFFASX1 \regfile_reg[6][0]  ( .D(n392), .CLK(clk), .SETB(rst), .Q(
        \regfile[6][0] ) );
  DFFARX1 \regfile_reg[7][0]  ( .D(n391), .CLK(clk), .RSTB(rst), .Q(
        \regfile[7][0] ) );
  DFFASX1 \regfile_reg[8][0]  ( .D(n390), .CLK(clk), .SETB(rst), .Q(
        \regfile[8][0] ) );
  DFFARX1 \regfile_reg[9][0]  ( .D(n389), .CLK(clk), .RSTB(rst), .Q(
        \regfile[9][0] ) );
  DFFASX1 \regfile_reg[10][0]  ( .D(n388), .CLK(clk), .SETB(rst), .Q(
        \regfile[10][0] ) );
  DFFARX1 \regfile_reg[11][0]  ( .D(n387), .CLK(clk), .RSTB(rst), .Q(
        \regfile[11][0] ) );
  DFFASX1 \regfile_reg[12][0]  ( .D(n386), .CLK(clk), .SETB(rst), .Q(
        \regfile[12][0] ) );
  DFFARX1 \regfile_reg[13][0]  ( .D(n385), .CLK(clk), .RSTB(rst), .Q(
        \regfile[13][0] ) );
  DFFASX1 \regfile_reg[14][0]  ( .D(n384), .CLK(clk), .SETB(rst), .Q(
        \regfile[14][0] ) );
  DFFARX1 \regfile_reg[15][0]  ( .D(n383), .CLK(clk), .RSTB(rst), .Q(
        \regfile[15][0] ) );
  pipealu_DW01_addsub_0 r308 ( .A({1'b0, IFID_A}), .B({1'b0, IFID_B}), .CI(
        1'b0), .ADD_SUB(n1494), .SUM({N255, N254, N253, N252, N251, N250, N249, 
        N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, 
        N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, 
        N224, N223}) );
  OR2X1 U895 ( .IN1(n1456), .IN2(n1002), .Q(n1004) );
  INVX0 U896 ( .INP(n1004), .ZN(n1008) );
  INVX0 U897 ( .INP(n1004), .ZN(n1009) );
  INVX0 U898 ( .INP(n1004), .ZN(n1010) );
  INVX0 U899 ( .INP(n1004), .ZN(n1011) );
  NOR2X1 U900 ( .IN1(n1001), .IN2(n1457), .QN(n1494) );
  MUX41X1 U901 ( .IN1(\regfile[12][0] ), .IN3(\regfile[14][0] ), .IN2(
        \regfile[13][0] ), .IN4(\regfile[15][0] ), .S0(N16), .S1(N15), .Q(
        n1012) );
  MUX41X1 U902 ( .IN1(\regfile[8][0] ), .IN3(\regfile[10][0] ), .IN2(
        \regfile[9][0] ), .IN4(\regfile[11][0] ), .S0(N16), .S1(N15), .Q(n1013) );
  MUX41X1 U903 ( .IN1(\regfile[4][0] ), .IN3(\regfile[6][0] ), .IN2(
        \regfile[5][0] ), .IN4(\regfile[7][0] ), .S0(N16), .S1(N15), .Q(n1014)
         );
  MUX41X1 U904 ( .IN1(\regfile[0][0] ), .IN3(\regfile[2][0] ), .IN2(
        \regfile[1][0] ), .IN4(\regfile[3][0] ), .S0(N16), .S1(N15), .Q(n1015)
         );
  MUX41X1 U905 ( .IN1(n1015), .IN3(n1013), .IN2(n1014), .IN4(n1012), .S0(N18), 
        .S1(N17), .Q(N55) );
  MUX41X1 U906 ( .IN1(\regfile[12][1] ), .IN3(\regfile[14][1] ), .IN2(
        \regfile[13][1] ), .IN4(\regfile[15][1] ), .S0(N16), .S1(N15), .Q(
        n1016) );
  MUX41X1 U907 ( .IN1(\regfile[8][1] ), .IN3(\regfile[10][1] ), .IN2(
        \regfile[9][1] ), .IN4(\regfile[11][1] ), .S0(N16), .S1(N15), .Q(n1017) );
  MUX41X1 U908 ( .IN1(\regfile[4][1] ), .IN3(\regfile[6][1] ), .IN2(
        \regfile[5][1] ), .IN4(\regfile[7][1] ), .S0(N16), .S1(N15), .Q(n1018)
         );
  MUX41X1 U909 ( .IN1(\regfile[0][1] ), .IN3(\regfile[2][1] ), .IN2(
        \regfile[1][1] ), .IN4(\regfile[3][1] ), .S0(N16), .S1(N15), .Q(n1019)
         );
  MUX41X1 U910 ( .IN1(n1019), .IN3(n1017), .IN2(n1018), .IN4(n1016), .S0(N18), 
        .S1(N17), .Q(N54) );
  MUX41X1 U911 ( .IN1(\regfile[12][2] ), .IN3(\regfile[14][2] ), .IN2(
        \regfile[13][2] ), .IN4(\regfile[15][2] ), .S0(N16), .S1(N15), .Q(
        n1020) );
  MUX41X1 U912 ( .IN1(\regfile[8][2] ), .IN3(\regfile[10][2] ), .IN2(
        \regfile[9][2] ), .IN4(\regfile[11][2] ), .S0(N16), .S1(N15), .Q(n1021) );
  MUX41X1 U913 ( .IN1(\regfile[4][2] ), .IN3(\regfile[6][2] ), .IN2(
        \regfile[5][2] ), .IN4(\regfile[7][2] ), .S0(N16), .S1(N15), .Q(n1022)
         );
  MUX41X1 U914 ( .IN1(\regfile[0][2] ), .IN3(\regfile[2][2] ), .IN2(
        \regfile[1][2] ), .IN4(\regfile[3][2] ), .S0(N16), .S1(N15), .Q(n1023)
         );
  MUX41X1 U915 ( .IN1(n1023), .IN3(n1021), .IN2(n1022), .IN4(n1020), .S0(N18), 
        .S1(N17), .Q(N53) );
  MUX41X1 U916 ( .IN1(\regfile[12][3] ), .IN3(\regfile[14][3] ), .IN2(
        \regfile[13][3] ), .IN4(\regfile[15][3] ), .S0(N16), .S1(N15), .Q(
        n1024) );
  MUX41X1 U917 ( .IN1(\regfile[8][3] ), .IN3(\regfile[10][3] ), .IN2(
        \regfile[9][3] ), .IN4(\regfile[11][3] ), .S0(N16), .S1(N15), .Q(n1025) );
  MUX41X1 U918 ( .IN1(\regfile[4][3] ), .IN3(\regfile[6][3] ), .IN2(
        \regfile[5][3] ), .IN4(\regfile[7][3] ), .S0(N16), .S1(N15), .Q(n1026)
         );
  MUX41X1 U919 ( .IN1(\regfile[0][3] ), .IN3(\regfile[2][3] ), .IN2(
        \regfile[1][3] ), .IN4(\regfile[3][3] ), .S0(N16), .S1(N15), .Q(n1027)
         );
  MUX41X1 U920 ( .IN1(n1027), .IN3(n1025), .IN2(n1026), .IN4(n1024), .S0(N18), 
        .S1(N17), .Q(N52) );
  MUX41X1 U921 ( .IN1(\regfile[12][4] ), .IN3(\regfile[14][4] ), .IN2(
        \regfile[13][4] ), .IN4(\regfile[15][4] ), .S0(N16), .S1(N15), .Q(
        n1028) );
  MUX41X1 U922 ( .IN1(\regfile[8][4] ), .IN3(\regfile[10][4] ), .IN2(
        \regfile[9][4] ), .IN4(\regfile[11][4] ), .S0(N16), .S1(N15), .Q(n1029) );
  MUX41X1 U923 ( .IN1(\regfile[4][4] ), .IN3(\regfile[6][4] ), .IN2(
        \regfile[5][4] ), .IN4(\regfile[7][4] ), .S0(N16), .S1(N15), .Q(n1030)
         );
  MUX41X1 U924 ( .IN1(\regfile[0][4] ), .IN3(\regfile[2][4] ), .IN2(
        \regfile[1][4] ), .IN4(\regfile[3][4] ), .S0(N16), .S1(N15), .Q(n1031)
         );
  MUX41X1 U925 ( .IN1(n1031), .IN3(n1029), .IN2(n1030), .IN4(n1028), .S0(N18), 
        .S1(N17), .Q(N51) );
  MUX41X1 U926 ( .IN1(\regfile[12][5] ), .IN3(\regfile[14][5] ), .IN2(
        \regfile[13][5] ), .IN4(\regfile[15][5] ), .S0(N16), .S1(N15), .Q(
        n1032) );
  MUX41X1 U927 ( .IN1(\regfile[8][5] ), .IN3(\regfile[10][5] ), .IN2(
        \regfile[9][5] ), .IN4(\regfile[11][5] ), .S0(N16), .S1(N15), .Q(n1033) );
  MUX41X1 U928 ( .IN1(\regfile[4][5] ), .IN3(\regfile[6][5] ), .IN2(
        \regfile[5][5] ), .IN4(\regfile[7][5] ), .S0(N16), .S1(N15), .Q(n1034)
         );
  MUX41X1 U929 ( .IN1(\regfile[0][5] ), .IN3(\regfile[2][5] ), .IN2(
        \regfile[1][5] ), .IN4(\regfile[3][5] ), .S0(N16), .S1(N15), .Q(n1035)
         );
  MUX41X1 U930 ( .IN1(n1035), .IN3(n1033), .IN2(n1034), .IN4(n1032), .S0(N18), 
        .S1(N17), .Q(N50) );
  MUX41X1 U931 ( .IN1(\regfile[12][6] ), .IN3(\regfile[14][6] ), .IN2(
        \regfile[13][6] ), .IN4(\regfile[15][6] ), .S0(N16), .S1(N15), .Q(
        n1036) );
  MUX41X1 U932 ( .IN1(\regfile[8][6] ), .IN3(\regfile[10][6] ), .IN2(
        \regfile[9][6] ), .IN4(\regfile[11][6] ), .S0(N16), .S1(N15), .Q(n1037) );
  MUX41X1 U933 ( .IN1(\regfile[4][6] ), .IN3(\regfile[6][6] ), .IN2(
        \regfile[5][6] ), .IN4(\regfile[7][6] ), .S0(N16), .S1(N15), .Q(n1038)
         );
  MUX41X1 U934 ( .IN1(\regfile[0][6] ), .IN3(\regfile[2][6] ), .IN2(
        \regfile[1][6] ), .IN4(\regfile[3][6] ), .S0(N16), .S1(N15), .Q(n1039)
         );
  MUX41X1 U935 ( .IN1(n1039), .IN3(n1037), .IN2(n1038), .IN4(n1036), .S0(N18), 
        .S1(N17), .Q(N49) );
  MUX41X1 U936 ( .IN1(\regfile[12][7] ), .IN3(\regfile[14][7] ), .IN2(
        \regfile[13][7] ), .IN4(\regfile[15][7] ), .S0(N16), .S1(N15), .Q(
        n1040) );
  MUX41X1 U937 ( .IN1(\regfile[8][7] ), .IN3(\regfile[10][7] ), .IN2(
        \regfile[9][7] ), .IN4(\regfile[11][7] ), .S0(N16), .S1(N15), .Q(n1041) );
  MUX41X1 U938 ( .IN1(\regfile[4][7] ), .IN3(\regfile[6][7] ), .IN2(
        \regfile[5][7] ), .IN4(\regfile[7][7] ), .S0(N16), .S1(N15), .Q(n1042)
         );
  MUX41X1 U939 ( .IN1(\regfile[0][7] ), .IN3(\regfile[2][7] ), .IN2(
        \regfile[1][7] ), .IN4(\regfile[3][7] ), .S0(N16), .S1(N15), .Q(n1043)
         );
  MUX41X1 U940 ( .IN1(n1043), .IN3(n1041), .IN2(n1042), .IN4(n1040), .S0(N18), 
        .S1(N17), .Q(N48) );
  MUX41X1 U941 ( .IN1(\regfile[12][8] ), .IN3(\regfile[14][8] ), .IN2(
        \regfile[13][8] ), .IN4(\regfile[15][8] ), .S0(N16), .S1(N15), .Q(
        n1044) );
  MUX41X1 U942 ( .IN1(\regfile[8][8] ), .IN3(\regfile[10][8] ), .IN2(
        \regfile[9][8] ), .IN4(\regfile[11][8] ), .S0(N16), .S1(N15), .Q(n1045) );
  MUX41X1 U943 ( .IN1(\regfile[4][8] ), .IN3(\regfile[6][8] ), .IN2(
        \regfile[5][8] ), .IN4(\regfile[7][8] ), .S0(N16), .S1(N15), .Q(n1046)
         );
  MUX41X1 U944 ( .IN1(\regfile[0][8] ), .IN3(\regfile[2][8] ), .IN2(
        \regfile[1][8] ), .IN4(\regfile[3][8] ), .S0(N16), .S1(N15), .Q(n1047)
         );
  MUX41X1 U945 ( .IN1(n1047), .IN3(n1045), .IN2(n1046), .IN4(n1044), .S0(N18), 
        .S1(N17), .Q(N47) );
  MUX41X1 U946 ( .IN1(\regfile[12][9] ), .IN3(\regfile[14][9] ), .IN2(
        \regfile[13][9] ), .IN4(\regfile[15][9] ), .S0(N16), .S1(N15), .Q(
        n1048) );
  MUX41X1 U947 ( .IN1(\regfile[8][9] ), .IN3(\regfile[10][9] ), .IN2(
        \regfile[9][9] ), .IN4(\regfile[11][9] ), .S0(N16), .S1(N15), .Q(n1049) );
  MUX41X1 U948 ( .IN1(\regfile[4][9] ), .IN3(\regfile[6][9] ), .IN2(
        \regfile[5][9] ), .IN4(\regfile[7][9] ), .S0(N16), .S1(N15), .Q(n1050)
         );
  MUX41X1 U949 ( .IN1(\regfile[0][9] ), .IN3(\regfile[2][9] ), .IN2(
        \regfile[1][9] ), .IN4(\regfile[3][9] ), .S0(N16), .S1(N15), .Q(n1051)
         );
  MUX41X1 U950 ( .IN1(n1051), .IN3(n1049), .IN2(n1050), .IN4(n1048), .S0(N18), 
        .S1(N17), .Q(N46) );
  MUX41X1 U951 ( .IN1(\regfile[12][10] ), .IN3(\regfile[14][10] ), .IN2(
        \regfile[13][10] ), .IN4(\regfile[15][10] ), .S0(N16), .S1(N15), .Q(
        n1052) );
  MUX41X1 U952 ( .IN1(\regfile[8][10] ), .IN3(\regfile[10][10] ), .IN2(
        \regfile[9][10] ), .IN4(\regfile[11][10] ), .S0(N16), .S1(N15), .Q(
        n1053) );
  MUX41X1 U953 ( .IN1(\regfile[4][10] ), .IN3(\regfile[6][10] ), .IN2(
        \regfile[5][10] ), .IN4(\regfile[7][10] ), .S0(N16), .S1(N15), .Q(
        n1054) );
  MUX41X1 U954 ( .IN1(\regfile[0][10] ), .IN3(\regfile[2][10] ), .IN2(
        \regfile[1][10] ), .IN4(\regfile[3][10] ), .S0(N16), .S1(N15), .Q(
        n1055) );
  MUX41X1 U955 ( .IN1(n1055), .IN3(n1053), .IN2(n1054), .IN4(n1052), .S0(N18), 
        .S1(N17), .Q(N45) );
  MUX41X1 U956 ( .IN1(\regfile[12][11] ), .IN3(\regfile[14][11] ), .IN2(
        \regfile[13][11] ), .IN4(\regfile[15][11] ), .S0(N16), .S1(N15), .Q(
        n1056) );
  MUX41X1 U957 ( .IN1(\regfile[8][11] ), .IN3(\regfile[10][11] ), .IN2(
        \regfile[9][11] ), .IN4(\regfile[11][11] ), .S0(N16), .S1(N15), .Q(
        n1057) );
  MUX41X1 U958 ( .IN1(\regfile[4][11] ), .IN3(\regfile[6][11] ), .IN2(
        \regfile[5][11] ), .IN4(\regfile[7][11] ), .S0(N16), .S1(N15), .Q(
        n1058) );
  MUX41X1 U959 ( .IN1(\regfile[0][11] ), .IN3(\regfile[2][11] ), .IN2(
        \regfile[1][11] ), .IN4(\regfile[3][11] ), .S0(N16), .S1(N15), .Q(
        n1059) );
  MUX41X1 U960 ( .IN1(n1059), .IN3(n1057), .IN2(n1058), .IN4(n1056), .S0(N18), 
        .S1(N17), .Q(N44) );
  MUX41X1 U961 ( .IN1(\regfile[12][12] ), .IN3(\regfile[14][12] ), .IN2(
        \regfile[13][12] ), .IN4(\regfile[15][12] ), .S0(N16), .S1(N15), .Q(
        n1060) );
  MUX41X1 U962 ( .IN1(\regfile[8][12] ), .IN3(\regfile[10][12] ), .IN2(
        \regfile[9][12] ), .IN4(\regfile[11][12] ), .S0(N16), .S1(N15), .Q(
        n1061) );
  MUX41X1 U963 ( .IN1(\regfile[4][12] ), .IN3(\regfile[6][12] ), .IN2(
        \regfile[5][12] ), .IN4(\regfile[7][12] ), .S0(N16), .S1(N15), .Q(
        n1062) );
  MUX41X1 U964 ( .IN1(\regfile[0][12] ), .IN3(\regfile[2][12] ), .IN2(
        \regfile[1][12] ), .IN4(\regfile[3][12] ), .S0(N16), .S1(N15), .Q(
        n1063) );
  MUX41X1 U965 ( .IN1(n1063), .IN3(n1061), .IN2(n1062), .IN4(n1060), .S0(N18), 
        .S1(N17), .Q(N43) );
  MUX41X1 U966 ( .IN1(\regfile[12][13] ), .IN3(\regfile[14][13] ), .IN2(
        \regfile[13][13] ), .IN4(\regfile[15][13] ), .S0(N16), .S1(N15), .Q(
        n1064) );
  MUX41X1 U967 ( .IN1(\regfile[8][13] ), .IN3(\regfile[10][13] ), .IN2(
        \regfile[9][13] ), .IN4(\regfile[11][13] ), .S0(N16), .S1(N15), .Q(
        n1065) );
  MUX41X1 U968 ( .IN1(\regfile[4][13] ), .IN3(\regfile[6][13] ), .IN2(
        \regfile[5][13] ), .IN4(\regfile[7][13] ), .S0(N16), .S1(N15), .Q(
        n1066) );
  MUX41X1 U969 ( .IN1(\regfile[0][13] ), .IN3(\regfile[2][13] ), .IN2(
        \regfile[1][13] ), .IN4(\regfile[3][13] ), .S0(N16), .S1(N15), .Q(
        n1067) );
  MUX41X1 U970 ( .IN1(n1067), .IN3(n1065), .IN2(n1066), .IN4(n1064), .S0(N18), 
        .S1(N17), .Q(N42) );
  MUX41X1 U971 ( .IN1(\regfile[12][14] ), .IN3(\regfile[14][14] ), .IN2(
        \regfile[13][14] ), .IN4(\regfile[15][14] ), .S0(N16), .S1(N15), .Q(
        n1068) );
  MUX41X1 U972 ( .IN1(\regfile[8][14] ), .IN3(\regfile[10][14] ), .IN2(
        \regfile[9][14] ), .IN4(\regfile[11][14] ), .S0(N16), .S1(N15), .Q(
        n1069) );
  MUX41X1 U973 ( .IN1(\regfile[4][14] ), .IN3(\regfile[6][14] ), .IN2(
        \regfile[5][14] ), .IN4(\regfile[7][14] ), .S0(N16), .S1(N15), .Q(
        n1070) );
  MUX41X1 U974 ( .IN1(\regfile[0][14] ), .IN3(\regfile[2][14] ), .IN2(
        \regfile[1][14] ), .IN4(\regfile[3][14] ), .S0(N16), .S1(N15), .Q(
        n1071) );
  MUX41X1 U975 ( .IN1(n1071), .IN3(n1069), .IN2(n1070), .IN4(n1068), .S0(N18), 
        .S1(N17), .Q(N41) );
  MUX41X1 U976 ( .IN1(\regfile[12][15] ), .IN3(\regfile[14][15] ), .IN2(
        \regfile[13][15] ), .IN4(\regfile[15][15] ), .S0(N16), .S1(N15), .Q(
        n1072) );
  MUX41X1 U977 ( .IN1(\regfile[8][15] ), .IN3(\regfile[10][15] ), .IN2(
        \regfile[9][15] ), .IN4(\regfile[11][15] ), .S0(N16), .S1(N15), .Q(
        n1073) );
  MUX41X1 U978 ( .IN1(\regfile[4][15] ), .IN3(\regfile[6][15] ), .IN2(
        \regfile[5][15] ), .IN4(\regfile[7][15] ), .S0(N16), .S1(N15), .Q(
        n1074) );
  MUX41X1 U979 ( .IN1(\regfile[0][15] ), .IN3(\regfile[2][15] ), .IN2(
        \regfile[1][15] ), .IN4(\regfile[3][15] ), .S0(N16), .S1(N15), .Q(
        n1075) );
  MUX41X1 U980 ( .IN1(n1075), .IN3(n1073), .IN2(n1074), .IN4(n1072), .S0(N18), 
        .S1(N17), .Q(N40) );
  MUX41X1 U981 ( .IN1(\regfile[12][16] ), .IN3(\regfile[14][16] ), .IN2(
        \regfile[13][16] ), .IN4(\regfile[15][16] ), .S0(N16), .S1(N15), .Q(
        n1076) );
  MUX41X1 U982 ( .IN1(\regfile[8][16] ), .IN3(\regfile[10][16] ), .IN2(
        \regfile[9][16] ), .IN4(\regfile[11][16] ), .S0(N16), .S1(N15), .Q(
        n1077) );
  MUX41X1 U983 ( .IN1(\regfile[4][16] ), .IN3(\regfile[6][16] ), .IN2(
        \regfile[5][16] ), .IN4(\regfile[7][16] ), .S0(N16), .S1(N15), .Q(
        n1078) );
  MUX41X1 U984 ( .IN1(\regfile[0][16] ), .IN3(\regfile[2][16] ), .IN2(
        \regfile[1][16] ), .IN4(\regfile[3][16] ), .S0(N16), .S1(N15), .Q(
        n1079) );
  MUX41X1 U985 ( .IN1(n1079), .IN3(n1077), .IN2(n1078), .IN4(n1076), .S0(N18), 
        .S1(N17), .Q(N39) );
  MUX41X1 U986 ( .IN1(\regfile[12][17] ), .IN3(\regfile[14][17] ), .IN2(
        \regfile[13][17] ), .IN4(\regfile[15][17] ), .S0(N16), .S1(N15), .Q(
        n1080) );
  MUX41X1 U987 ( .IN1(\regfile[8][17] ), .IN3(\regfile[10][17] ), .IN2(
        \regfile[9][17] ), .IN4(\regfile[11][17] ), .S0(N16), .S1(N15), .Q(
        n1081) );
  MUX41X1 U988 ( .IN1(\regfile[4][17] ), .IN3(\regfile[6][17] ), .IN2(
        \regfile[5][17] ), .IN4(\regfile[7][17] ), .S0(N16), .S1(N15), .Q(
        n1082) );
  MUX41X1 U989 ( .IN1(\regfile[0][17] ), .IN3(\regfile[2][17] ), .IN2(
        \regfile[1][17] ), .IN4(\regfile[3][17] ), .S0(N16), .S1(N15), .Q(
        n1083) );
  MUX41X1 U990 ( .IN1(n1083), .IN3(n1081), .IN2(n1082), .IN4(n1080), .S0(N18), 
        .S1(N17), .Q(N38) );
  MUX41X1 U991 ( .IN1(\regfile[12][18] ), .IN3(\regfile[14][18] ), .IN2(
        \regfile[13][18] ), .IN4(\regfile[15][18] ), .S0(N16), .S1(N15), .Q(
        n1084) );
  MUX41X1 U992 ( .IN1(\regfile[8][18] ), .IN3(\regfile[10][18] ), .IN2(
        \regfile[9][18] ), .IN4(\regfile[11][18] ), .S0(N16), .S1(N15), .Q(
        n1085) );
  MUX41X1 U993 ( .IN1(\regfile[4][18] ), .IN3(\regfile[6][18] ), .IN2(
        \regfile[5][18] ), .IN4(\regfile[7][18] ), .S0(N16), .S1(N15), .Q(
        n1086) );
  MUX41X1 U994 ( .IN1(\regfile[0][18] ), .IN3(\regfile[2][18] ), .IN2(
        \regfile[1][18] ), .IN4(\regfile[3][18] ), .S0(N16), .S1(N15), .Q(
        n1087) );
  MUX41X1 U995 ( .IN1(n1087), .IN3(n1085), .IN2(n1086), .IN4(n1084), .S0(N18), 
        .S1(N17), .Q(N37) );
  MUX41X1 U996 ( .IN1(\regfile[12][19] ), .IN3(\regfile[14][19] ), .IN2(
        \regfile[13][19] ), .IN4(\regfile[15][19] ), .S0(N16), .S1(N15), .Q(
        n1088) );
  MUX41X1 U997 ( .IN1(\regfile[8][19] ), .IN3(\regfile[10][19] ), .IN2(
        \regfile[9][19] ), .IN4(\regfile[11][19] ), .S0(N16), .S1(N15), .Q(
        n1089) );
  MUX41X1 U998 ( .IN1(\regfile[4][19] ), .IN3(\regfile[6][19] ), .IN2(
        \regfile[5][19] ), .IN4(\regfile[7][19] ), .S0(N16), .S1(N15), .Q(
        n1090) );
  MUX41X1 U999 ( .IN1(\regfile[0][19] ), .IN3(\regfile[2][19] ), .IN2(
        \regfile[1][19] ), .IN4(\regfile[3][19] ), .S0(N16), .S1(N15), .Q(
        n1091) );
  MUX41X1 U1000 ( .IN1(n1091), .IN3(n1089), .IN2(n1090), .IN4(n1088), .S0(N18), 
        .S1(N17), .Q(N36) );
  MUX41X1 U1001 ( .IN1(\regfile[12][20] ), .IN3(\regfile[14][20] ), .IN2(
        \regfile[13][20] ), .IN4(\regfile[15][20] ), .S0(N16), .S1(N15), .Q(
        n1092) );
  MUX41X1 U1002 ( .IN1(\regfile[8][20] ), .IN3(\regfile[10][20] ), .IN2(
        \regfile[9][20] ), .IN4(\regfile[11][20] ), .S0(N16), .S1(N15), .Q(
        n1093) );
  MUX41X1 U1003 ( .IN1(\regfile[4][20] ), .IN3(\regfile[6][20] ), .IN2(
        \regfile[5][20] ), .IN4(\regfile[7][20] ), .S0(N16), .S1(N15), .Q(
        n1094) );
  MUX41X1 U1004 ( .IN1(\regfile[0][20] ), .IN3(\regfile[2][20] ), .IN2(
        \regfile[1][20] ), .IN4(\regfile[3][20] ), .S0(N16), .S1(N15), .Q(
        n1095) );
  MUX41X1 U1005 ( .IN1(n1095), .IN3(n1093), .IN2(n1094), .IN4(n1092), .S0(N18), 
        .S1(N17), .Q(N35) );
  MUX41X1 U1006 ( .IN1(\regfile[12][21] ), .IN3(\regfile[14][21] ), .IN2(
        \regfile[13][21] ), .IN4(\regfile[15][21] ), .S0(N16), .S1(N15), .Q(
        n1096) );
  MUX41X1 U1007 ( .IN1(\regfile[8][21] ), .IN3(\regfile[10][21] ), .IN2(
        \regfile[9][21] ), .IN4(\regfile[11][21] ), .S0(N16), .S1(N15), .Q(
        n1097) );
  MUX41X1 U1008 ( .IN1(\regfile[4][21] ), .IN3(\regfile[6][21] ), .IN2(
        \regfile[5][21] ), .IN4(\regfile[7][21] ), .S0(N16), .S1(N15), .Q(
        n1098) );
  MUX41X1 U1009 ( .IN1(\regfile[0][21] ), .IN3(\regfile[2][21] ), .IN2(
        \regfile[1][21] ), .IN4(\regfile[3][21] ), .S0(N16), .S1(N15), .Q(
        n1099) );
  MUX41X1 U1010 ( .IN1(n1099), .IN3(n1097), .IN2(n1098), .IN4(n1096), .S0(N18), 
        .S1(N17), .Q(N34) );
  MUX41X1 U1011 ( .IN1(\regfile[12][22] ), .IN3(\regfile[14][22] ), .IN2(
        \regfile[13][22] ), .IN4(\regfile[15][22] ), .S0(N16), .S1(N15), .Q(
        n1100) );
  MUX41X1 U1012 ( .IN1(\regfile[8][22] ), .IN3(\regfile[10][22] ), .IN2(
        \regfile[9][22] ), .IN4(\regfile[11][22] ), .S0(N16), .S1(N15), .Q(
        n1101) );
  MUX41X1 U1013 ( .IN1(\regfile[4][22] ), .IN3(\regfile[6][22] ), .IN2(
        \regfile[5][22] ), .IN4(\regfile[7][22] ), .S0(N16), .S1(N15), .Q(
        n1102) );
  MUX41X1 U1014 ( .IN1(\regfile[0][22] ), .IN3(\regfile[2][22] ), .IN2(
        \regfile[1][22] ), .IN4(\regfile[3][22] ), .S0(N16), .S1(N15), .Q(
        n1103) );
  MUX41X1 U1015 ( .IN1(n1103), .IN3(n1101), .IN2(n1102), .IN4(n1100), .S0(N18), 
        .S1(N17), .Q(N33) );
  MUX41X1 U1016 ( .IN1(\regfile[12][23] ), .IN3(\regfile[14][23] ), .IN2(
        \regfile[13][23] ), .IN4(\regfile[15][23] ), .S0(N16), .S1(N15), .Q(
        n1104) );
  MUX41X1 U1017 ( .IN1(\regfile[8][23] ), .IN3(\regfile[10][23] ), .IN2(
        \regfile[9][23] ), .IN4(\regfile[11][23] ), .S0(N16), .S1(N15), .Q(
        n1105) );
  MUX41X1 U1018 ( .IN1(\regfile[4][23] ), .IN3(\regfile[6][23] ), .IN2(
        \regfile[5][23] ), .IN4(\regfile[7][23] ), .S0(N16), .S1(N15), .Q(
        n1106) );
  MUX41X1 U1019 ( .IN1(\regfile[0][23] ), .IN3(\regfile[2][23] ), .IN2(
        \regfile[1][23] ), .IN4(\regfile[3][23] ), .S0(N16), .S1(N15), .Q(
        n1107) );
  MUX41X1 U1020 ( .IN1(n1107), .IN3(n1105), .IN2(n1106), .IN4(n1104), .S0(N18), 
        .S1(N17), .Q(N32) );
  MUX41X1 U1021 ( .IN1(\regfile[12][24] ), .IN3(\regfile[14][24] ), .IN2(
        \regfile[13][24] ), .IN4(\regfile[15][24] ), .S0(N16), .S1(N15), .Q(
        n1108) );
  MUX41X1 U1022 ( .IN1(\regfile[8][24] ), .IN3(\regfile[10][24] ), .IN2(
        \regfile[9][24] ), .IN4(\regfile[11][24] ), .S0(N16), .S1(N15), .Q(
        n1109) );
  MUX41X1 U1023 ( .IN1(\regfile[4][24] ), .IN3(\regfile[6][24] ), .IN2(
        \regfile[5][24] ), .IN4(\regfile[7][24] ), .S0(N16), .S1(N15), .Q(
        n1110) );
  MUX41X1 U1024 ( .IN1(\regfile[0][24] ), .IN3(\regfile[2][24] ), .IN2(
        \regfile[1][24] ), .IN4(\regfile[3][24] ), .S0(N16), .S1(N15), .Q(
        n1111) );
  MUX41X1 U1025 ( .IN1(n1111), .IN3(n1109), .IN2(n1110), .IN4(n1108), .S0(N18), 
        .S1(N17), .Q(N31) );
  MUX41X1 U1026 ( .IN1(\regfile[12][25] ), .IN3(\regfile[14][25] ), .IN2(
        \regfile[13][25] ), .IN4(\regfile[15][25] ), .S0(N16), .S1(N15), .Q(
        n1112) );
  MUX41X1 U1027 ( .IN1(\regfile[8][25] ), .IN3(\regfile[10][25] ), .IN2(
        \regfile[9][25] ), .IN4(\regfile[11][25] ), .S0(N16), .S1(N15), .Q(
        n1113) );
  MUX41X1 U1028 ( .IN1(\regfile[4][25] ), .IN3(\regfile[6][25] ), .IN2(
        \regfile[5][25] ), .IN4(\regfile[7][25] ), .S0(N16), .S1(N15), .Q(
        n1114) );
  MUX41X1 U1029 ( .IN1(\regfile[0][25] ), .IN3(\regfile[2][25] ), .IN2(
        \regfile[1][25] ), .IN4(\regfile[3][25] ), .S0(N16), .S1(N15), .Q(
        n1115) );
  MUX41X1 U1030 ( .IN1(n1115), .IN3(n1113), .IN2(n1114), .IN4(n1112), .S0(N18), 
        .S1(N17), .Q(N30) );
  MUX41X1 U1031 ( .IN1(\regfile[12][26] ), .IN3(\regfile[14][26] ), .IN2(
        \regfile[13][26] ), .IN4(\regfile[15][26] ), .S0(N16), .S1(N15), .Q(
        n1116) );
  MUX41X1 U1032 ( .IN1(\regfile[8][26] ), .IN3(\regfile[10][26] ), .IN2(
        \regfile[9][26] ), .IN4(\regfile[11][26] ), .S0(N16), .S1(N15), .Q(
        n1117) );
  MUX41X1 U1033 ( .IN1(\regfile[4][26] ), .IN3(\regfile[6][26] ), .IN2(
        \regfile[5][26] ), .IN4(\regfile[7][26] ), .S0(N16), .S1(N15), .Q(
        n1118) );
  MUX41X1 U1034 ( .IN1(\regfile[0][26] ), .IN3(\regfile[2][26] ), .IN2(
        \regfile[1][26] ), .IN4(\regfile[3][26] ), .S0(N16), .S1(N15), .Q(
        n1119) );
  MUX41X1 U1035 ( .IN1(n1119), .IN3(n1117), .IN2(n1118), .IN4(n1116), .S0(N18), 
        .S1(N17), .Q(N29) );
  MUX41X1 U1036 ( .IN1(\regfile[12][27] ), .IN3(\regfile[14][27] ), .IN2(
        \regfile[13][27] ), .IN4(\regfile[15][27] ), .S0(N16), .S1(N15), .Q(
        n1120) );
  MUX41X1 U1037 ( .IN1(\regfile[8][27] ), .IN3(\regfile[10][27] ), .IN2(
        \regfile[9][27] ), .IN4(\regfile[11][27] ), .S0(N16), .S1(N15), .Q(
        n1121) );
  MUX41X1 U1038 ( .IN1(\regfile[4][27] ), .IN3(\regfile[6][27] ), .IN2(
        \regfile[5][27] ), .IN4(\regfile[7][27] ), .S0(N16), .S1(N15), .Q(
        n1122) );
  MUX41X1 U1039 ( .IN1(\regfile[0][27] ), .IN3(\regfile[2][27] ), .IN2(
        \regfile[1][27] ), .IN4(\regfile[3][27] ), .S0(N16), .S1(N15), .Q(
        n1123) );
  MUX41X1 U1040 ( .IN1(n1123), .IN3(n1121), .IN2(n1122), .IN4(n1120), .S0(N18), 
        .S1(N17), .Q(N28) );
  MUX41X1 U1041 ( .IN1(\regfile[12][28] ), .IN3(\regfile[14][28] ), .IN2(
        \regfile[13][28] ), .IN4(\regfile[15][28] ), .S0(N16), .S1(N15), .Q(
        n1124) );
  MUX41X1 U1042 ( .IN1(\regfile[8][28] ), .IN3(\regfile[10][28] ), .IN2(
        \regfile[9][28] ), .IN4(\regfile[11][28] ), .S0(N16), .S1(N15), .Q(
        n1125) );
  MUX41X1 U1043 ( .IN1(\regfile[4][28] ), .IN3(\regfile[6][28] ), .IN2(
        \regfile[5][28] ), .IN4(\regfile[7][28] ), .S0(N16), .S1(N15), .Q(
        n1126) );
  MUX41X1 U1044 ( .IN1(\regfile[0][28] ), .IN3(\regfile[2][28] ), .IN2(
        \regfile[1][28] ), .IN4(\regfile[3][28] ), .S0(N16), .S1(N15), .Q(
        n1127) );
  MUX41X1 U1045 ( .IN1(n1127), .IN3(n1125), .IN2(n1126), .IN4(n1124), .S0(N18), 
        .S1(N17), .Q(N27) );
  MUX41X1 U1046 ( .IN1(\regfile[12][29] ), .IN3(\regfile[14][29] ), .IN2(
        \regfile[13][29] ), .IN4(\regfile[15][29] ), .S0(N16), .S1(N15), .Q(
        n1128) );
  MUX41X1 U1047 ( .IN1(\regfile[8][29] ), .IN3(\regfile[10][29] ), .IN2(
        \regfile[9][29] ), .IN4(\regfile[11][29] ), .S0(N16), .S1(N15), .Q(
        n1129) );
  MUX41X1 U1048 ( .IN1(\regfile[4][29] ), .IN3(\regfile[6][29] ), .IN2(
        \regfile[5][29] ), .IN4(\regfile[7][29] ), .S0(N16), .S1(N15), .Q(
        n1130) );
  MUX41X1 U1049 ( .IN1(\regfile[0][29] ), .IN3(\regfile[2][29] ), .IN2(
        \regfile[1][29] ), .IN4(\regfile[3][29] ), .S0(N16), .S1(N15), .Q(
        n1131) );
  MUX41X1 U1050 ( .IN1(n1131), .IN3(n1129), .IN2(n1130), .IN4(n1128), .S0(N18), 
        .S1(N17), .Q(N26) );
  MUX41X1 U1051 ( .IN1(\regfile[12][30] ), .IN3(\regfile[14][30] ), .IN2(
        \regfile[13][30] ), .IN4(\regfile[15][30] ), .S0(N16), .S1(N15), .Q(
        n1132) );
  MUX41X1 U1052 ( .IN1(\regfile[8][30] ), .IN3(\regfile[10][30] ), .IN2(
        \regfile[9][30] ), .IN4(\regfile[11][30] ), .S0(N16), .S1(N15), .Q(
        n1133) );
  MUX41X1 U1053 ( .IN1(\regfile[4][30] ), .IN3(\regfile[6][30] ), .IN2(
        \regfile[5][30] ), .IN4(\regfile[7][30] ), .S0(N16), .S1(N15), .Q(
        n1134) );
  MUX41X1 U1054 ( .IN1(\regfile[0][30] ), .IN3(\regfile[2][30] ), .IN2(
        \regfile[1][30] ), .IN4(\regfile[3][30] ), .S0(N16), .S1(N15), .Q(
        n1135) );
  MUX41X1 U1055 ( .IN1(n1135), .IN3(n1133), .IN2(n1134), .IN4(n1132), .S0(N18), 
        .S1(N17), .Q(N25) );
  MUX41X1 U1056 ( .IN1(\regfile[12][31] ), .IN3(\regfile[14][31] ), .IN2(
        \regfile[13][31] ), .IN4(\regfile[15][31] ), .S0(N16), .S1(N15), .Q(
        n1136) );
  MUX41X1 U1057 ( .IN1(\regfile[8][31] ), .IN3(\regfile[10][31] ), .IN2(
        \regfile[9][31] ), .IN4(\regfile[11][31] ), .S0(N16), .S1(N15), .Q(
        n1137) );
  MUX41X1 U1058 ( .IN1(\regfile[4][31] ), .IN3(\regfile[6][31] ), .IN2(
        \regfile[5][31] ), .IN4(\regfile[7][31] ), .S0(N16), .S1(N15), .Q(
        n1138) );
  MUX41X1 U1059 ( .IN1(\regfile[0][31] ), .IN3(\regfile[2][31] ), .IN2(
        \regfile[1][31] ), .IN4(\regfile[3][31] ), .S0(N16), .S1(N15), .Q(
        n1139) );
  MUX41X1 U1060 ( .IN1(n1139), .IN3(n1137), .IN2(n1138), .IN4(n1136), .S0(N18), 
        .S1(N17), .Q(N24) );
  MUX41X1 U1061 ( .IN1(\regfile[12][0] ), .IN3(\regfile[14][0] ), .IN2(
        \regfile[13][0] ), .IN4(\regfile[15][0] ), .S0(N20), .S1(N19), .Q(
        n1140) );
  MUX41X1 U1062 ( .IN1(\regfile[8][0] ), .IN3(\regfile[10][0] ), .IN2(
        \regfile[9][0] ), .IN4(\regfile[11][0] ), .S0(N20), .S1(N19), .Q(n1141) );
  MUX41X1 U1063 ( .IN1(\regfile[4][0] ), .IN3(\regfile[6][0] ), .IN2(
        \regfile[5][0] ), .IN4(\regfile[7][0] ), .S0(N20), .S1(N19), .Q(n1142)
         );
  MUX41X1 U1064 ( .IN1(\regfile[0][0] ), .IN3(\regfile[2][0] ), .IN2(
        \regfile[1][0] ), .IN4(\regfile[3][0] ), .S0(N20), .S1(N19), .Q(n1143)
         );
  MUX41X1 U1065 ( .IN1(n1143), .IN3(n1141), .IN2(n1142), .IN4(n1140), .S0(N22), 
        .S1(N21), .Q(N87) );
  MUX41X1 U1066 ( .IN1(\regfile[12][1] ), .IN3(\regfile[14][1] ), .IN2(
        \regfile[13][1] ), .IN4(\regfile[15][1] ), .S0(N20), .S1(N19), .Q(
        n1144) );
  MUX41X1 U1067 ( .IN1(\regfile[8][1] ), .IN3(\regfile[10][1] ), .IN2(
        \regfile[9][1] ), .IN4(\regfile[11][1] ), .S0(N20), .S1(N19), .Q(n1145) );
  MUX41X1 U1068 ( .IN1(\regfile[4][1] ), .IN3(\regfile[6][1] ), .IN2(
        \regfile[5][1] ), .IN4(\regfile[7][1] ), .S0(N20), .S1(N19), .Q(n1146)
         );
  MUX41X1 U1069 ( .IN1(\regfile[0][1] ), .IN3(\regfile[2][1] ), .IN2(
        \regfile[1][1] ), .IN4(\regfile[3][1] ), .S0(N20), .S1(N19), .Q(n1147)
         );
  MUX41X1 U1070 ( .IN1(n1147), .IN3(n1145), .IN2(n1146), .IN4(n1144), .S0(N22), 
        .S1(N21), .Q(N86) );
  MUX41X1 U1071 ( .IN1(\regfile[12][2] ), .IN3(\regfile[14][2] ), .IN2(
        \regfile[13][2] ), .IN4(\regfile[15][2] ), .S0(N20), .S1(N19), .Q(
        n1148) );
  MUX41X1 U1072 ( .IN1(\regfile[8][2] ), .IN3(\regfile[10][2] ), .IN2(
        \regfile[9][2] ), .IN4(\regfile[11][2] ), .S0(N20), .S1(N19), .Q(n1149) );
  MUX41X1 U1073 ( .IN1(\regfile[4][2] ), .IN3(\regfile[6][2] ), .IN2(
        \regfile[5][2] ), .IN4(\regfile[7][2] ), .S0(N20), .S1(N19), .Q(n1150)
         );
  MUX41X1 U1074 ( .IN1(\regfile[0][2] ), .IN3(\regfile[2][2] ), .IN2(
        \regfile[1][2] ), .IN4(\regfile[3][2] ), .S0(N20), .S1(N19), .Q(n1151)
         );
  MUX41X1 U1075 ( .IN1(n1151), .IN3(n1149), .IN2(n1150), .IN4(n1148), .S0(N22), 
        .S1(N21), .Q(N85) );
  MUX41X1 U1076 ( .IN1(\regfile[12][3] ), .IN3(\regfile[14][3] ), .IN2(
        \regfile[13][3] ), .IN4(\regfile[15][3] ), .S0(N20), .S1(N19), .Q(
        n1152) );
  MUX41X1 U1077 ( .IN1(\regfile[8][3] ), .IN3(\regfile[10][3] ), .IN2(
        \regfile[9][3] ), .IN4(\regfile[11][3] ), .S0(N20), .S1(N19), .Q(n1153) );
  MUX41X1 U1078 ( .IN1(\regfile[4][3] ), .IN3(\regfile[6][3] ), .IN2(
        \regfile[5][3] ), .IN4(\regfile[7][3] ), .S0(N20), .S1(N19), .Q(n1154)
         );
  MUX41X1 U1079 ( .IN1(\regfile[0][3] ), .IN3(\regfile[2][3] ), .IN2(
        \regfile[1][3] ), .IN4(\regfile[3][3] ), .S0(N20), .S1(N19), .Q(n1155)
         );
  MUX41X1 U1080 ( .IN1(n1155), .IN3(n1153), .IN2(n1154), .IN4(n1152), .S0(N22), 
        .S1(N21), .Q(N84) );
  MUX41X1 U1081 ( .IN1(\regfile[12][4] ), .IN3(\regfile[14][4] ), .IN2(
        \regfile[13][4] ), .IN4(\regfile[15][4] ), .S0(N20), .S1(N19), .Q(
        n1156) );
  MUX41X1 U1082 ( .IN1(\regfile[8][4] ), .IN3(\regfile[10][4] ), .IN2(
        \regfile[9][4] ), .IN4(\regfile[11][4] ), .S0(N20), .S1(N19), .Q(n1157) );
  MUX41X1 U1083 ( .IN1(\regfile[4][4] ), .IN3(\regfile[6][4] ), .IN2(
        \regfile[5][4] ), .IN4(\regfile[7][4] ), .S0(N20), .S1(N19), .Q(n1158)
         );
  MUX41X1 U1084 ( .IN1(\regfile[0][4] ), .IN3(\regfile[2][4] ), .IN2(
        \regfile[1][4] ), .IN4(\regfile[3][4] ), .S0(N20), .S1(N19), .Q(n1159)
         );
  MUX41X1 U1085 ( .IN1(n1159), .IN3(n1157), .IN2(n1158), .IN4(n1156), .S0(N22), 
        .S1(N21), .Q(N83) );
  MUX41X1 U1086 ( .IN1(\regfile[12][5] ), .IN3(\regfile[14][5] ), .IN2(
        \regfile[13][5] ), .IN4(\regfile[15][5] ), .S0(N20), .S1(N19), .Q(
        n1160) );
  MUX41X1 U1087 ( .IN1(\regfile[8][5] ), .IN3(\regfile[10][5] ), .IN2(
        \regfile[9][5] ), .IN4(\regfile[11][5] ), .S0(N20), .S1(N19), .Q(n1161) );
  MUX41X1 U1088 ( .IN1(\regfile[4][5] ), .IN3(\regfile[6][5] ), .IN2(
        \regfile[5][5] ), .IN4(\regfile[7][5] ), .S0(N20), .S1(N19), .Q(n1162)
         );
  MUX41X1 U1089 ( .IN1(\regfile[0][5] ), .IN3(\regfile[2][5] ), .IN2(
        \regfile[1][5] ), .IN4(\regfile[3][5] ), .S0(N20), .S1(N19), .Q(n1163)
         );
  MUX41X1 U1090 ( .IN1(n1163), .IN3(n1161), .IN2(n1162), .IN4(n1160), .S0(N22), 
        .S1(N21), .Q(N82) );
  MUX41X1 U1091 ( .IN1(\regfile[12][6] ), .IN3(\regfile[14][6] ), .IN2(
        \regfile[13][6] ), .IN4(\regfile[15][6] ), .S0(N20), .S1(N19), .Q(
        n1164) );
  MUX41X1 U1092 ( .IN1(\regfile[8][6] ), .IN3(\regfile[10][6] ), .IN2(
        \regfile[9][6] ), .IN4(\regfile[11][6] ), .S0(N20), .S1(N19), .Q(n1165) );
  MUX41X1 U1093 ( .IN1(\regfile[4][6] ), .IN3(\regfile[6][6] ), .IN2(
        \regfile[5][6] ), .IN4(\regfile[7][6] ), .S0(N20), .S1(N19), .Q(n1166)
         );
  MUX41X1 U1094 ( .IN1(\regfile[0][6] ), .IN3(\regfile[2][6] ), .IN2(
        \regfile[1][6] ), .IN4(\regfile[3][6] ), .S0(N20), .S1(N19), .Q(n1167)
         );
  MUX41X1 U1095 ( .IN1(n1167), .IN3(n1165), .IN2(n1166), .IN4(n1164), .S0(N22), 
        .S1(N21), .Q(N81) );
  MUX41X1 U1096 ( .IN1(\regfile[12][7] ), .IN3(\regfile[14][7] ), .IN2(
        \regfile[13][7] ), .IN4(\regfile[15][7] ), .S0(N20), .S1(N19), .Q(
        n1168) );
  MUX41X1 U1097 ( .IN1(\regfile[8][7] ), .IN3(\regfile[10][7] ), .IN2(
        \regfile[9][7] ), .IN4(\regfile[11][7] ), .S0(N20), .S1(N19), .Q(n1169) );
  MUX41X1 U1098 ( .IN1(\regfile[4][7] ), .IN3(\regfile[6][7] ), .IN2(
        \regfile[5][7] ), .IN4(\regfile[7][7] ), .S0(N20), .S1(N19), .Q(n1170)
         );
  MUX41X1 U1099 ( .IN1(\regfile[0][7] ), .IN3(\regfile[2][7] ), .IN2(
        \regfile[1][7] ), .IN4(\regfile[3][7] ), .S0(N20), .S1(N19), .Q(n1171)
         );
  MUX41X1 U1100 ( .IN1(n1171), .IN3(n1169), .IN2(n1170), .IN4(n1168), .S0(N22), 
        .S1(N21), .Q(N80) );
  MUX41X1 U1101 ( .IN1(\regfile[12][8] ), .IN3(\regfile[14][8] ), .IN2(
        \regfile[13][8] ), .IN4(\regfile[15][8] ), .S0(N20), .S1(N19), .Q(
        n1172) );
  MUX41X1 U1102 ( .IN1(\regfile[8][8] ), .IN3(\regfile[10][8] ), .IN2(
        \regfile[9][8] ), .IN4(\regfile[11][8] ), .S0(N20), .S1(N19), .Q(n1173) );
  MUX41X1 U1103 ( .IN1(\regfile[4][8] ), .IN3(\regfile[6][8] ), .IN2(
        \regfile[5][8] ), .IN4(\regfile[7][8] ), .S0(N20), .S1(N19), .Q(n1174)
         );
  MUX41X1 U1104 ( .IN1(\regfile[0][8] ), .IN3(\regfile[2][8] ), .IN2(
        \regfile[1][8] ), .IN4(\regfile[3][8] ), .S0(N20), .S1(N19), .Q(n1175)
         );
  MUX41X1 U1105 ( .IN1(n1175), .IN3(n1173), .IN2(n1174), .IN4(n1172), .S0(N22), 
        .S1(N21), .Q(N79) );
  MUX41X1 U1106 ( .IN1(\regfile[12][9] ), .IN3(\regfile[14][9] ), .IN2(
        \regfile[13][9] ), .IN4(\regfile[15][9] ), .S0(N20), .S1(N19), .Q(
        n1176) );
  MUX41X1 U1107 ( .IN1(\regfile[8][9] ), .IN3(\regfile[10][9] ), .IN2(
        \regfile[9][9] ), .IN4(\regfile[11][9] ), .S0(N20), .S1(N19), .Q(n1177) );
  MUX41X1 U1108 ( .IN1(\regfile[4][9] ), .IN3(\regfile[6][9] ), .IN2(
        \regfile[5][9] ), .IN4(\regfile[7][9] ), .S0(N20), .S1(N19), .Q(n1178)
         );
  MUX41X1 U1109 ( .IN1(\regfile[0][9] ), .IN3(\regfile[2][9] ), .IN2(
        \regfile[1][9] ), .IN4(\regfile[3][9] ), .S0(N20), .S1(N19), .Q(n1179)
         );
  MUX41X1 U1110 ( .IN1(n1179), .IN3(n1177), .IN2(n1178), .IN4(n1176), .S0(N22), 
        .S1(N21), .Q(N78) );
  MUX41X1 U1111 ( .IN1(\regfile[12][10] ), .IN3(\regfile[14][10] ), .IN2(
        \regfile[13][10] ), .IN4(\regfile[15][10] ), .S0(N20), .S1(N19), .Q(
        n1180) );
  MUX41X1 U1112 ( .IN1(\regfile[8][10] ), .IN3(\regfile[10][10] ), .IN2(
        \regfile[9][10] ), .IN4(\regfile[11][10] ), .S0(N20), .S1(N19), .Q(
        n1181) );
  MUX41X1 U1113 ( .IN1(\regfile[4][10] ), .IN3(\regfile[6][10] ), .IN2(
        \regfile[5][10] ), .IN4(\regfile[7][10] ), .S0(N20), .S1(N19), .Q(
        n1182) );
  MUX41X1 U1114 ( .IN1(\regfile[0][10] ), .IN3(\regfile[2][10] ), .IN2(
        \regfile[1][10] ), .IN4(\regfile[3][10] ), .S0(N20), .S1(N19), .Q(
        n1183) );
  MUX41X1 U1115 ( .IN1(n1183), .IN3(n1181), .IN2(n1182), .IN4(n1180), .S0(N22), 
        .S1(N21), .Q(N77) );
  MUX41X1 U1116 ( .IN1(\regfile[12][11] ), .IN3(\regfile[14][11] ), .IN2(
        \regfile[13][11] ), .IN4(\regfile[15][11] ), .S0(N20), .S1(N19), .Q(
        n1184) );
  MUX41X1 U1117 ( .IN1(\regfile[8][11] ), .IN3(\regfile[10][11] ), .IN2(
        \regfile[9][11] ), .IN4(\regfile[11][11] ), .S0(N20), .S1(N19), .Q(
        n1185) );
  MUX41X1 U1118 ( .IN1(\regfile[4][11] ), .IN3(\regfile[6][11] ), .IN2(
        \regfile[5][11] ), .IN4(\regfile[7][11] ), .S0(N20), .S1(N19), .Q(
        n1186) );
  MUX41X1 U1119 ( .IN1(\regfile[0][11] ), .IN3(\regfile[2][11] ), .IN2(
        \regfile[1][11] ), .IN4(\regfile[3][11] ), .S0(N20), .S1(N19), .Q(
        n1187) );
  MUX41X1 U1120 ( .IN1(n1187), .IN3(n1185), .IN2(n1186), .IN4(n1184), .S0(N22), 
        .S1(N21), .Q(N76) );
  MUX41X1 U1121 ( .IN1(\regfile[12][12] ), .IN3(\regfile[14][12] ), .IN2(
        \regfile[13][12] ), .IN4(\regfile[15][12] ), .S0(N20), .S1(N19), .Q(
        n1188) );
  MUX41X1 U1122 ( .IN1(\regfile[8][12] ), .IN3(\regfile[10][12] ), .IN2(
        \regfile[9][12] ), .IN4(\regfile[11][12] ), .S0(N20), .S1(N19), .Q(
        n1189) );
  MUX41X1 U1123 ( .IN1(\regfile[4][12] ), .IN3(\regfile[6][12] ), .IN2(
        \regfile[5][12] ), .IN4(\regfile[7][12] ), .S0(N20), .S1(N19), .Q(
        n1190) );
  MUX41X1 U1124 ( .IN1(\regfile[0][12] ), .IN3(\regfile[2][12] ), .IN2(
        \regfile[1][12] ), .IN4(\regfile[3][12] ), .S0(N20), .S1(N19), .Q(
        n1191) );
  MUX41X1 U1125 ( .IN1(n1191), .IN3(n1189), .IN2(n1190), .IN4(n1188), .S0(N22), 
        .S1(N21), .Q(N75) );
  MUX41X1 U1126 ( .IN1(\regfile[12][13] ), .IN3(\regfile[14][13] ), .IN2(
        \regfile[13][13] ), .IN4(\regfile[15][13] ), .S0(N20), .S1(N19), .Q(
        n1192) );
  MUX41X1 U1127 ( .IN1(\regfile[8][13] ), .IN3(\regfile[10][13] ), .IN2(
        \regfile[9][13] ), .IN4(\regfile[11][13] ), .S0(N20), .S1(N19), .Q(
        n1193) );
  MUX41X1 U1128 ( .IN1(\regfile[4][13] ), .IN3(\regfile[6][13] ), .IN2(
        \regfile[5][13] ), .IN4(\regfile[7][13] ), .S0(N20), .S1(N19), .Q(
        n1194) );
  MUX41X1 U1129 ( .IN1(\regfile[0][13] ), .IN3(\regfile[2][13] ), .IN2(
        \regfile[1][13] ), .IN4(\regfile[3][13] ), .S0(N20), .S1(N19), .Q(
        n1195) );
  MUX41X1 U1130 ( .IN1(n1195), .IN3(n1193), .IN2(n1194), .IN4(n1192), .S0(N22), 
        .S1(N21), .Q(N74) );
  MUX41X1 U1131 ( .IN1(\regfile[12][14] ), .IN3(\regfile[14][14] ), .IN2(
        \regfile[13][14] ), .IN4(\regfile[15][14] ), .S0(N20), .S1(N19), .Q(
        n1196) );
  MUX41X1 U1132 ( .IN1(\regfile[8][14] ), .IN3(\regfile[10][14] ), .IN2(
        \regfile[9][14] ), .IN4(\regfile[11][14] ), .S0(N20), .S1(N19), .Q(
        n1197) );
  MUX41X1 U1133 ( .IN1(\regfile[4][14] ), .IN3(\regfile[6][14] ), .IN2(
        \regfile[5][14] ), .IN4(\regfile[7][14] ), .S0(N20), .S1(N19), .Q(
        n1198) );
  MUX41X1 U1134 ( .IN1(\regfile[0][14] ), .IN3(\regfile[2][14] ), .IN2(
        \regfile[1][14] ), .IN4(\regfile[3][14] ), .S0(N20), .S1(N19), .Q(
        n1199) );
  MUX41X1 U1135 ( .IN1(n1199), .IN3(n1197), .IN2(n1198), .IN4(n1196), .S0(N22), 
        .S1(N21), .Q(N73) );
  MUX41X1 U1136 ( .IN1(\regfile[12][15] ), .IN3(\regfile[14][15] ), .IN2(
        \regfile[13][15] ), .IN4(\regfile[15][15] ), .S0(N20), .S1(N19), .Q(
        n1200) );
  MUX41X1 U1137 ( .IN1(\regfile[8][15] ), .IN3(\regfile[10][15] ), .IN2(
        \regfile[9][15] ), .IN4(\regfile[11][15] ), .S0(N20), .S1(N19), .Q(
        n1201) );
  MUX41X1 U1138 ( .IN1(\regfile[4][15] ), .IN3(\regfile[6][15] ), .IN2(
        \regfile[5][15] ), .IN4(\regfile[7][15] ), .S0(N20), .S1(N19), .Q(
        n1202) );
  MUX41X1 U1139 ( .IN1(\regfile[0][15] ), .IN3(\regfile[2][15] ), .IN2(
        \regfile[1][15] ), .IN4(\regfile[3][15] ), .S0(N20), .S1(N19), .Q(
        n1203) );
  MUX41X1 U1140 ( .IN1(n1203), .IN3(n1201), .IN2(n1202), .IN4(n1200), .S0(N22), 
        .S1(N21), .Q(N72) );
  MUX41X1 U1141 ( .IN1(\regfile[12][16] ), .IN3(\regfile[14][16] ), .IN2(
        \regfile[13][16] ), .IN4(\regfile[15][16] ), .S0(N20), .S1(N19), .Q(
        n1204) );
  MUX41X1 U1142 ( .IN1(\regfile[8][16] ), .IN3(\regfile[10][16] ), .IN2(
        \regfile[9][16] ), .IN4(\regfile[11][16] ), .S0(N20), .S1(N19), .Q(
        n1205) );
  MUX41X1 U1143 ( .IN1(\regfile[4][16] ), .IN3(\regfile[6][16] ), .IN2(
        \regfile[5][16] ), .IN4(\regfile[7][16] ), .S0(N20), .S1(N19), .Q(
        n1206) );
  MUX41X1 U1144 ( .IN1(\regfile[0][16] ), .IN3(\regfile[2][16] ), .IN2(
        \regfile[1][16] ), .IN4(\regfile[3][16] ), .S0(N20), .S1(N19), .Q(
        n1207) );
  MUX41X1 U1145 ( .IN1(n1207), .IN3(n1205), .IN2(n1206), .IN4(n1204), .S0(N22), 
        .S1(N21), .Q(N71) );
  MUX41X1 U1146 ( .IN1(\regfile[12][17] ), .IN3(\regfile[14][17] ), .IN2(
        \regfile[13][17] ), .IN4(\regfile[15][17] ), .S0(N20), .S1(N19), .Q(
        n1208) );
  MUX41X1 U1147 ( .IN1(\regfile[8][17] ), .IN3(\regfile[10][17] ), .IN2(
        \regfile[9][17] ), .IN4(\regfile[11][17] ), .S0(N20), .S1(N19), .Q(
        n1209) );
  MUX41X1 U1148 ( .IN1(\regfile[4][17] ), .IN3(\regfile[6][17] ), .IN2(
        \regfile[5][17] ), .IN4(\regfile[7][17] ), .S0(N20), .S1(N19), .Q(
        n1210) );
  MUX41X1 U1149 ( .IN1(\regfile[0][17] ), .IN3(\regfile[2][17] ), .IN2(
        \regfile[1][17] ), .IN4(\regfile[3][17] ), .S0(N20), .S1(N19), .Q(
        n1211) );
  MUX41X1 U1150 ( .IN1(n1211), .IN3(n1209), .IN2(n1210), .IN4(n1208), .S0(N22), 
        .S1(N21), .Q(N70) );
  MUX41X1 U1151 ( .IN1(\regfile[12][18] ), .IN3(\regfile[14][18] ), .IN2(
        \regfile[13][18] ), .IN4(\regfile[15][18] ), .S0(N20), .S1(N19), .Q(
        n1212) );
  MUX41X1 U1152 ( .IN1(\regfile[8][18] ), .IN3(\regfile[10][18] ), .IN2(
        \regfile[9][18] ), .IN4(\regfile[11][18] ), .S0(N20), .S1(N19), .Q(
        n1213) );
  MUX41X1 U1153 ( .IN1(\regfile[4][18] ), .IN3(\regfile[6][18] ), .IN2(
        \regfile[5][18] ), .IN4(\regfile[7][18] ), .S0(N20), .S1(N19), .Q(
        n1214) );
  MUX41X1 U1154 ( .IN1(\regfile[0][18] ), .IN3(\regfile[2][18] ), .IN2(
        \regfile[1][18] ), .IN4(\regfile[3][18] ), .S0(N20), .S1(N19), .Q(
        n1215) );
  MUX41X1 U1155 ( .IN1(n1215), .IN3(n1213), .IN2(n1214), .IN4(n1212), .S0(N22), 
        .S1(N21), .Q(N69) );
  MUX41X1 U1156 ( .IN1(\regfile[12][19] ), .IN3(\regfile[14][19] ), .IN2(
        \regfile[13][19] ), .IN4(\regfile[15][19] ), .S0(N20), .S1(N19), .Q(
        n1216) );
  MUX41X1 U1157 ( .IN1(\regfile[8][19] ), .IN3(\regfile[10][19] ), .IN2(
        \regfile[9][19] ), .IN4(\regfile[11][19] ), .S0(N20), .S1(N19), .Q(
        n1217) );
  MUX41X1 U1158 ( .IN1(\regfile[4][19] ), .IN3(\regfile[6][19] ), .IN2(
        \regfile[5][19] ), .IN4(\regfile[7][19] ), .S0(N20), .S1(N19), .Q(
        n1218) );
  MUX41X1 U1159 ( .IN1(\regfile[0][19] ), .IN3(\regfile[2][19] ), .IN2(
        \regfile[1][19] ), .IN4(\regfile[3][19] ), .S0(N20), .S1(N19), .Q(
        n1219) );
  MUX41X1 U1160 ( .IN1(n1219), .IN3(n1217), .IN2(n1218), .IN4(n1216), .S0(N22), 
        .S1(N21), .Q(N68) );
  MUX41X1 U1161 ( .IN1(\regfile[12][20] ), .IN3(\regfile[14][20] ), .IN2(
        \regfile[13][20] ), .IN4(\regfile[15][20] ), .S0(N20), .S1(N19), .Q(
        n1220) );
  MUX41X1 U1162 ( .IN1(\regfile[8][20] ), .IN3(\regfile[10][20] ), .IN2(
        \regfile[9][20] ), .IN4(\regfile[11][20] ), .S0(N20), .S1(N19), .Q(
        n1221) );
  MUX41X1 U1163 ( .IN1(\regfile[4][20] ), .IN3(\regfile[6][20] ), .IN2(
        \regfile[5][20] ), .IN4(\regfile[7][20] ), .S0(N20), .S1(N19), .Q(
        n1222) );
  MUX41X1 U1164 ( .IN1(\regfile[0][20] ), .IN3(\regfile[2][20] ), .IN2(
        \regfile[1][20] ), .IN4(\regfile[3][20] ), .S0(N20), .S1(N19), .Q(
        n1223) );
  MUX41X1 U1165 ( .IN1(n1223), .IN3(n1221), .IN2(n1222), .IN4(n1220), .S0(N22), 
        .S1(N21), .Q(N67) );
  MUX41X1 U1166 ( .IN1(\regfile[12][21] ), .IN3(\regfile[14][21] ), .IN2(
        \regfile[13][21] ), .IN4(\regfile[15][21] ), .S0(N20), .S1(N19), .Q(
        n1224) );
  MUX41X1 U1167 ( .IN1(\regfile[8][21] ), .IN3(\regfile[10][21] ), .IN2(
        \regfile[9][21] ), .IN4(\regfile[11][21] ), .S0(N20), .S1(N19), .Q(
        n1225) );
  MUX41X1 U1168 ( .IN1(\regfile[4][21] ), .IN3(\regfile[6][21] ), .IN2(
        \regfile[5][21] ), .IN4(\regfile[7][21] ), .S0(N20), .S1(N19), .Q(
        n1226) );
  MUX41X1 U1169 ( .IN1(\regfile[0][21] ), .IN3(\regfile[2][21] ), .IN2(
        \regfile[1][21] ), .IN4(\regfile[3][21] ), .S0(N20), .S1(N19), .Q(
        n1227) );
  MUX41X1 U1170 ( .IN1(n1227), .IN3(n1225), .IN2(n1226), .IN4(n1224), .S0(N22), 
        .S1(N21), .Q(N66) );
  MUX41X1 U1171 ( .IN1(\regfile[12][22] ), .IN3(\regfile[14][22] ), .IN2(
        \regfile[13][22] ), .IN4(\regfile[15][22] ), .S0(N20), .S1(N19), .Q(
        n1228) );
  MUX41X1 U1172 ( .IN1(\regfile[8][22] ), .IN3(\regfile[10][22] ), .IN2(
        \regfile[9][22] ), .IN4(\regfile[11][22] ), .S0(N20), .S1(N19), .Q(
        n1229) );
  MUX41X1 U1173 ( .IN1(\regfile[4][22] ), .IN3(\regfile[6][22] ), .IN2(
        \regfile[5][22] ), .IN4(\regfile[7][22] ), .S0(N20), .S1(N19), .Q(
        n1230) );
  MUX41X1 U1174 ( .IN1(\regfile[0][22] ), .IN3(\regfile[2][22] ), .IN2(
        \regfile[1][22] ), .IN4(\regfile[3][22] ), .S0(N20), .S1(N19), .Q(
        n1231) );
  MUX41X1 U1175 ( .IN1(n1231), .IN3(n1229), .IN2(n1230), .IN4(n1228), .S0(N22), 
        .S1(N21), .Q(N65) );
  MUX41X1 U1176 ( .IN1(\regfile[12][23] ), .IN3(\regfile[14][23] ), .IN2(
        \regfile[13][23] ), .IN4(\regfile[15][23] ), .S0(N20), .S1(N19), .Q(
        n1232) );
  MUX41X1 U1177 ( .IN1(\regfile[8][23] ), .IN3(\regfile[10][23] ), .IN2(
        \regfile[9][23] ), .IN4(\regfile[11][23] ), .S0(N20), .S1(N19), .Q(
        n1233) );
  MUX41X1 U1178 ( .IN1(\regfile[4][23] ), .IN3(\regfile[6][23] ), .IN2(
        \regfile[5][23] ), .IN4(\regfile[7][23] ), .S0(N20), .S1(N19), .Q(
        n1234) );
  MUX41X1 U1179 ( .IN1(\regfile[0][23] ), .IN3(\regfile[2][23] ), .IN2(
        \regfile[1][23] ), .IN4(\regfile[3][23] ), .S0(N20), .S1(N19), .Q(
        n1235) );
  MUX41X1 U1180 ( .IN1(n1235), .IN3(n1233), .IN2(n1234), .IN4(n1232), .S0(N22), 
        .S1(N21), .Q(N64) );
  MUX41X1 U1181 ( .IN1(\regfile[12][24] ), .IN3(\regfile[14][24] ), .IN2(
        \regfile[13][24] ), .IN4(\regfile[15][24] ), .S0(N20), .S1(N19), .Q(
        n1236) );
  MUX41X1 U1182 ( .IN1(\regfile[8][24] ), .IN3(\regfile[10][24] ), .IN2(
        \regfile[9][24] ), .IN4(\regfile[11][24] ), .S0(N20), .S1(N19), .Q(
        n1237) );
  MUX41X1 U1183 ( .IN1(\regfile[4][24] ), .IN3(\regfile[6][24] ), .IN2(
        \regfile[5][24] ), .IN4(\regfile[7][24] ), .S0(N20), .S1(N19), .Q(
        n1238) );
  MUX41X1 U1184 ( .IN1(\regfile[0][24] ), .IN3(\regfile[2][24] ), .IN2(
        \regfile[1][24] ), .IN4(\regfile[3][24] ), .S0(N20), .S1(N19), .Q(
        n1239) );
  MUX41X1 U1185 ( .IN1(n1239), .IN3(n1237), .IN2(n1238), .IN4(n1236), .S0(N22), 
        .S1(N21), .Q(N63) );
  MUX41X1 U1186 ( .IN1(\regfile[12][25] ), .IN3(\regfile[14][25] ), .IN2(
        \regfile[13][25] ), .IN4(\regfile[15][25] ), .S0(N20), .S1(N19), .Q(
        n1240) );
  MUX41X1 U1187 ( .IN1(\regfile[8][25] ), .IN3(\regfile[10][25] ), .IN2(
        \regfile[9][25] ), .IN4(\regfile[11][25] ), .S0(N20), .S1(N19), .Q(
        n1241) );
  MUX41X1 U1188 ( .IN1(\regfile[4][25] ), .IN3(\regfile[6][25] ), .IN2(
        \regfile[5][25] ), .IN4(\regfile[7][25] ), .S0(N20), .S1(N19), .Q(
        n1242) );
  MUX41X1 U1189 ( .IN1(\regfile[0][25] ), .IN3(\regfile[2][25] ), .IN2(
        \regfile[1][25] ), .IN4(\regfile[3][25] ), .S0(N20), .S1(N19), .Q(
        n1243) );
  MUX41X1 U1190 ( .IN1(n1243), .IN3(n1241), .IN2(n1242), .IN4(n1240), .S0(N22), 
        .S1(N21), .Q(N62) );
  MUX41X1 U1191 ( .IN1(\regfile[12][26] ), .IN3(\regfile[14][26] ), .IN2(
        \regfile[13][26] ), .IN4(\regfile[15][26] ), .S0(N20), .S1(N19), .Q(
        n1244) );
  MUX41X1 U1192 ( .IN1(\regfile[8][26] ), .IN3(\regfile[10][26] ), .IN2(
        \regfile[9][26] ), .IN4(\regfile[11][26] ), .S0(N20), .S1(N19), .Q(
        n1245) );
  MUX41X1 U1193 ( .IN1(\regfile[4][26] ), .IN3(\regfile[6][26] ), .IN2(
        \regfile[5][26] ), .IN4(\regfile[7][26] ), .S0(N20), .S1(N19), .Q(
        n1246) );
  MUX41X1 U1194 ( .IN1(\regfile[0][26] ), .IN3(\regfile[2][26] ), .IN2(
        \regfile[1][26] ), .IN4(\regfile[3][26] ), .S0(N20), .S1(N19), .Q(
        n1247) );
  MUX41X1 U1195 ( .IN1(n1247), .IN3(n1245), .IN2(n1246), .IN4(n1244), .S0(N22), 
        .S1(N21), .Q(N61) );
  MUX41X1 U1196 ( .IN1(\regfile[12][27] ), .IN3(\regfile[14][27] ), .IN2(
        \regfile[13][27] ), .IN4(\regfile[15][27] ), .S0(N20), .S1(N19), .Q(
        n1248) );
  MUX41X1 U1197 ( .IN1(\regfile[8][27] ), .IN3(\regfile[10][27] ), .IN2(
        \regfile[9][27] ), .IN4(\regfile[11][27] ), .S0(N20), .S1(N19), .Q(
        n1249) );
  MUX41X1 U1198 ( .IN1(\regfile[4][27] ), .IN3(\regfile[6][27] ), .IN2(
        \regfile[5][27] ), .IN4(\regfile[7][27] ), .S0(N20), .S1(N19), .Q(
        n1250) );
  MUX41X1 U1199 ( .IN1(\regfile[0][27] ), .IN3(\regfile[2][27] ), .IN2(
        \regfile[1][27] ), .IN4(\regfile[3][27] ), .S0(N20), .S1(N19), .Q(
        n1251) );
  MUX41X1 U1200 ( .IN1(n1251), .IN3(n1249), .IN2(n1250), .IN4(n1248), .S0(N22), 
        .S1(N21), .Q(N60) );
  MUX41X1 U1201 ( .IN1(\regfile[12][28] ), .IN3(\regfile[14][28] ), .IN2(
        \regfile[13][28] ), .IN4(\regfile[15][28] ), .S0(N20), .S1(N19), .Q(
        n1252) );
  MUX41X1 U1202 ( .IN1(\regfile[8][28] ), .IN3(\regfile[10][28] ), .IN2(
        \regfile[9][28] ), .IN4(\regfile[11][28] ), .S0(N20), .S1(N19), .Q(
        n1253) );
  MUX41X1 U1203 ( .IN1(\regfile[4][28] ), .IN3(\regfile[6][28] ), .IN2(
        \regfile[5][28] ), .IN4(\regfile[7][28] ), .S0(N20), .S1(N19), .Q(
        n1254) );
  MUX41X1 U1204 ( .IN1(\regfile[0][28] ), .IN3(\regfile[2][28] ), .IN2(
        \regfile[1][28] ), .IN4(\regfile[3][28] ), .S0(N20), .S1(N19), .Q(
        n1255) );
  MUX41X1 U1205 ( .IN1(n1255), .IN3(n1253), .IN2(n1254), .IN4(n1252), .S0(N22), 
        .S1(N21), .Q(N59) );
  MUX41X1 U1206 ( .IN1(\regfile[12][29] ), .IN3(\regfile[14][29] ), .IN2(
        \regfile[13][29] ), .IN4(\regfile[15][29] ), .S0(N20), .S1(N19), .Q(
        n1256) );
  MUX41X1 U1207 ( .IN1(\regfile[8][29] ), .IN3(\regfile[10][29] ), .IN2(
        \regfile[9][29] ), .IN4(\regfile[11][29] ), .S0(N20), .S1(N19), .Q(
        n1257) );
  MUX41X1 U1208 ( .IN1(\regfile[4][29] ), .IN3(\regfile[6][29] ), .IN2(
        \regfile[5][29] ), .IN4(\regfile[7][29] ), .S0(N20), .S1(N19), .Q(
        n1258) );
  MUX41X1 U1209 ( .IN1(\regfile[0][29] ), .IN3(\regfile[2][29] ), .IN2(
        \regfile[1][29] ), .IN4(\regfile[3][29] ), .S0(N20), .S1(N19), .Q(
        n1259) );
  MUX41X1 U1210 ( .IN1(n1259), .IN3(n1257), .IN2(n1258), .IN4(n1256), .S0(N22), 
        .S1(N21), .Q(N58) );
  MUX41X1 U1211 ( .IN1(\regfile[12][30] ), .IN3(\regfile[14][30] ), .IN2(
        \regfile[13][30] ), .IN4(\regfile[15][30] ), .S0(N20), .S1(N19), .Q(
        n1260) );
  MUX41X1 U1212 ( .IN1(\regfile[8][30] ), .IN3(\regfile[10][30] ), .IN2(
        \regfile[9][30] ), .IN4(\regfile[11][30] ), .S0(N20), .S1(N19), .Q(
        n1261) );
  MUX41X1 U1213 ( .IN1(\regfile[4][30] ), .IN3(\regfile[6][30] ), .IN2(
        \regfile[5][30] ), .IN4(\regfile[7][30] ), .S0(N20), .S1(N19), .Q(
        n1262) );
  MUX41X1 U1214 ( .IN1(\regfile[0][30] ), .IN3(\regfile[2][30] ), .IN2(
        \regfile[1][30] ), .IN4(\regfile[3][30] ), .S0(N20), .S1(N19), .Q(
        n1263) );
  MUX41X1 U1215 ( .IN1(n1263), .IN3(n1261), .IN2(n1262), .IN4(n1260), .S0(N22), 
        .S1(N21), .Q(N57) );
  MUX41X1 U1216 ( .IN1(\regfile[12][31] ), .IN3(\regfile[14][31] ), .IN2(
        \regfile[13][31] ), .IN4(\regfile[15][31] ), .S0(N20), .S1(N19), .Q(
        n1264) );
  MUX41X1 U1217 ( .IN1(\regfile[8][31] ), .IN3(\regfile[10][31] ), .IN2(
        \regfile[9][31] ), .IN4(\regfile[11][31] ), .S0(N20), .S1(N19), .Q(
        n1265) );
  MUX41X1 U1218 ( .IN1(\regfile[4][31] ), .IN3(\regfile[6][31] ), .IN2(
        \regfile[5][31] ), .IN4(\regfile[7][31] ), .S0(N20), .S1(N19), .Q(
        n1266) );
  MUX41X1 U1219 ( .IN1(\regfile[0][31] ), .IN3(\regfile[2][31] ), .IN2(
        \regfile[1][31] ), .IN4(\regfile[3][31] ), .S0(N20), .S1(N19), .Q(
        n1267) );
  MUX41X1 U1220 ( .IN1(n1267), .IN3(n1265), .IN2(n1266), .IN4(n1264), .S0(N22), 
        .S1(N21), .Q(N56) );
  MUX21X1 U1221 ( .IN1(IFID_B[31]), .IN2(N56), .S(rst), .Q(n998) );
  MUX21X1 U1222 ( .IN1(IFID_B[30]), .IN2(N57), .S(rst), .Q(n997) );
  MUX21X1 U1223 ( .IN1(IFID_B[29]), .IN2(N58), .S(rst), .Q(n996) );
  MUX21X1 U1224 ( .IN1(IFID_B[28]), .IN2(N59), .S(rst), .Q(n995) );
  MUX21X1 U1225 ( .IN1(IFID_B[27]), .IN2(N60), .S(rst), .Q(n994) );
  MUX21X1 U1226 ( .IN1(IFID_B[26]), .IN2(N61), .S(rst), .Q(n993) );
  MUX21X1 U1227 ( .IN1(IFID_B[25]), .IN2(N62), .S(rst), .Q(n992) );
  MUX21X1 U1228 ( .IN1(IFID_B[24]), .IN2(N63), .S(rst), .Q(n991) );
  MUX21X1 U1229 ( .IN1(IFID_B[23]), .IN2(N64), .S(rst), .Q(n990) );
  MUX21X1 U1230 ( .IN1(IFID_B[22]), .IN2(N65), .S(rst), .Q(n989) );
  MUX21X1 U1231 ( .IN1(IFID_B[21]), .IN2(N66), .S(rst), .Q(n988) );
  MUX21X1 U1232 ( .IN1(IFID_B[20]), .IN2(N67), .S(rst), .Q(n987) );
  MUX21X1 U1233 ( .IN1(IFID_B[19]), .IN2(N68), .S(rst), .Q(n986) );
  MUX21X1 U1234 ( .IN1(IFID_B[18]), .IN2(N69), .S(rst), .Q(n985) );
  MUX21X1 U1235 ( .IN1(IFID_B[17]), .IN2(N70), .S(rst), .Q(n984) );
  MUX21X1 U1236 ( .IN1(IFID_B[16]), .IN2(N71), .S(rst), .Q(n983) );
  MUX21X1 U1237 ( .IN1(IFID_B[15]), .IN2(N72), .S(rst), .Q(n982) );
  MUX21X1 U1238 ( .IN1(IFID_B[14]), .IN2(N73), .S(rst), .Q(n981) );
  MUX21X1 U1239 ( .IN1(IFID_B[13]), .IN2(N74), .S(rst), .Q(n980) );
  MUX21X1 U1240 ( .IN1(IFID_B[12]), .IN2(N75), .S(rst), .Q(n979) );
  MUX21X1 U1241 ( .IN1(IFID_B[11]), .IN2(N76), .S(rst), .Q(n978) );
  MUX21X1 U1242 ( .IN1(IFID_B[10]), .IN2(N77), .S(rst), .Q(n977) );
  MUX21X1 U1243 ( .IN1(IFID_B[9]), .IN2(N78), .S(rst), .Q(n976) );
  MUX21X1 U1244 ( .IN1(IFID_B[8]), .IN2(N79), .S(rst), .Q(n975) );
  MUX21X1 U1245 ( .IN1(IFID_B[7]), .IN2(N80), .S(rst), .Q(n974) );
  MUX21X1 U1246 ( .IN1(IFID_B[6]), .IN2(N81), .S(rst), .Q(n973) );
  MUX21X1 U1247 ( .IN1(IFID_B[5]), .IN2(N82), .S(rst), .Q(n972) );
  MUX21X1 U1248 ( .IN1(IFID_B[4]), .IN2(N83), .S(rst), .Q(n971) );
  MUX21X1 U1249 ( .IN1(IFID_B[3]), .IN2(N84), .S(rst), .Q(n970) );
  MUX21X1 U1250 ( .IN1(IFID_B[2]), .IN2(N85), .S(rst), .Q(n969) );
  MUX21X1 U1251 ( .IN1(IFID_B[1]), .IN2(N86), .S(rst), .Q(n968) );
  MUX21X1 U1252 ( .IN1(IFID_B[0]), .IN2(N87), .S(rst), .Q(n967) );
  MUX21X1 U1253 ( .IN1(n1488), .IN2(instr[15]), .S(rst), .Q(n966) );
  MUX21X1 U1254 ( .IN1(n1487), .IN2(instr[14]), .S(rst), .Q(n965) );
  MUX21X1 U1255 ( .IN1(n1486), .IN2(instr[13]), .S(rst), .Q(n964) );
  MUX21X1 U1256 ( .IN1(n1485), .IN2(instr[12]), .S(rst), .Q(n963) );
  MUX21X1 U1257 ( .IN1(IFID_A[31]), .IN2(N24), .S(rst), .Q(n962) );
  MUX21X1 U1258 ( .IN1(IFID_A[30]), .IN2(N25), .S(rst), .Q(n961) );
  MUX21X1 U1259 ( .IN1(IFID_A[29]), .IN2(N26), .S(rst), .Q(n960) );
  MUX21X1 U1260 ( .IN1(IFID_A[28]), .IN2(N27), .S(rst), .Q(n959) );
  MUX21X1 U1261 ( .IN1(IFID_A[27]), .IN2(N28), .S(rst), .Q(n958) );
  MUX21X1 U1262 ( .IN1(IFID_A[26]), .IN2(N29), .S(rst), .Q(n957) );
  MUX21X1 U1263 ( .IN1(IFID_A[25]), .IN2(N30), .S(rst), .Q(n956) );
  MUX21X1 U1264 ( .IN1(IFID_A[24]), .IN2(N31), .S(rst), .Q(n955) );
  MUX21X1 U1265 ( .IN1(IFID_A[23]), .IN2(N32), .S(rst), .Q(n954) );
  MUX21X1 U1266 ( .IN1(IFID_A[22]), .IN2(N33), .S(rst), .Q(n953) );
  MUX21X1 U1267 ( .IN1(IFID_A[21]), .IN2(N34), .S(rst), .Q(n952) );
  MUX21X1 U1268 ( .IN1(IFID_A[20]), .IN2(N35), .S(rst), .Q(n951) );
  MUX21X1 U1269 ( .IN1(IFID_A[19]), .IN2(N36), .S(rst), .Q(n950) );
  MUX21X1 U1270 ( .IN1(IFID_A[18]), .IN2(N37), .S(rst), .Q(n949) );
  MUX21X1 U1271 ( .IN1(IFID_A[17]), .IN2(N38), .S(rst), .Q(n948) );
  MUX21X1 U1272 ( .IN1(IFID_A[16]), .IN2(N39), .S(rst), .Q(n947) );
  MUX21X1 U1273 ( .IN1(IFID_A[15]), .IN2(N40), .S(rst), .Q(n946) );
  MUX21X1 U1274 ( .IN1(IFID_A[14]), .IN2(N41), .S(rst), .Q(n945) );
  MUX21X1 U1275 ( .IN1(IFID_A[13]), .IN2(N42), .S(rst), .Q(n944) );
  MUX21X1 U1276 ( .IN1(IFID_A[12]), .IN2(N43), .S(rst), .Q(n943) );
  MUX21X1 U1277 ( .IN1(IFID_A[11]), .IN2(N44), .S(rst), .Q(n942) );
  MUX21X1 U1278 ( .IN1(IFID_A[10]), .IN2(N45), .S(rst), .Q(n941) );
  MUX21X1 U1279 ( .IN1(IFID_A[9]), .IN2(N46), .S(rst), .Q(n940) );
  MUX21X1 U1280 ( .IN1(IFID_A[8]), .IN2(N47), .S(rst), .Q(n939) );
  MUX21X1 U1281 ( .IN1(IFID_A[7]), .IN2(N48), .S(rst), .Q(n938) );
  MUX21X1 U1282 ( .IN1(IFID_A[6]), .IN2(N49), .S(rst), .Q(n937) );
  MUX21X1 U1283 ( .IN1(IFID_A[5]), .IN2(N50), .S(rst), .Q(n936) );
  MUX21X1 U1284 ( .IN1(IFID_A[4]), .IN2(N51), .S(rst), .Q(n935) );
  MUX21X1 U1285 ( .IN1(IFID_A[3]), .IN2(N52), .S(rst), .Q(n934) );
  MUX21X1 U1286 ( .IN1(IFID_A[2]), .IN2(N53), .S(rst), .Q(n933) );
  MUX21X1 U1287 ( .IN1(IFID_A[1]), .IN2(N54), .S(rst), .Q(n932) );
  MUX21X1 U1288 ( .IN1(IFID_A[0]), .IN2(N55), .S(rst), .Q(n931) );
  MUX21X1 U1289 ( .IN1(IFID_dest[3]), .IN2(instr[3]), .S(rst), .Q(n930) );
  MUX21X1 U1290 ( .IN1(IFID_dest[2]), .IN2(instr[2]), .S(rst), .Q(n929) );
  MUX21X1 U1291 ( .IN1(IFID_dest[1]), .IN2(instr[1]), .S(rst), .Q(n928) );
  MUX21X1 U1292 ( .IN1(IFID_dest[0]), .IN2(instr[0]), .S(rst), .Q(n927) );
  AO221X1 U1293 ( .IN1(n1268), .IN2(AluOut[31]), .IN3(N254), .IN4(n1269), 
        .IN5(n1270), .Q(n926) );
  AO21X1 U1294 ( .IN1(n1010), .IN2(IFID_A[31]), .IN3(n1271), .Q(n1270) );
  MUX21X1 U1295 ( .IN1(n1272), .IN2(n1273), .S(IFID_B[31]), .Q(n1271) );
  AO21X1 U1296 ( .IN1(n1274), .IN2(IFID_A[31]), .IN3(n1011), .Q(n1273) );
  NOR2X0 U1297 ( .IN1(n1275), .IN2(IFID_A[31]), .QN(n1272) );
  MUX21X1 U1298 ( .IN1(\regfile[0][31] ), .IN2(AluOut[31]), .S(n1276), .Q(n925) );
  MUX21X1 U1299 ( .IN1(\regfile[1][31] ), .IN2(AluOut[31]), .S(n1277), .Q(n924) );
  MUX21X1 U1300 ( .IN1(\regfile[2][31] ), .IN2(AluOut[31]), .S(n1278), .Q(n923) );
  MUX21X1 U1301 ( .IN1(\regfile[3][31] ), .IN2(AluOut[31]), .S(n1279), .Q(n922) );
  MUX21X1 U1302 ( .IN1(\regfile[4][31] ), .IN2(AluOut[31]), .S(n1280), .Q(n921) );
  MUX21X1 U1303 ( .IN1(\regfile[5][31] ), .IN2(AluOut[31]), .S(n1281), .Q(n920) );
  MUX21X1 U1304 ( .IN1(\regfile[6][31] ), .IN2(AluOut[31]), .S(n1282), .Q(n919) );
  MUX21X1 U1305 ( .IN1(\regfile[7][31] ), .IN2(AluOut[31]), .S(n1283), .Q(n918) );
  MUX21X1 U1306 ( .IN1(\regfile[8][31] ), .IN2(AluOut[31]), .S(n1284), .Q(n917) );
  MUX21X1 U1307 ( .IN1(\regfile[9][31] ), .IN2(AluOut[31]), .S(n1285), .Q(n916) );
  MUX21X1 U1308 ( .IN1(\regfile[10][31] ), .IN2(AluOut[31]), .S(n1286), .Q(
        n915) );
  MUX21X1 U1309 ( .IN1(\regfile[11][31] ), .IN2(AluOut[31]), .S(n1287), .Q(
        n914) );
  MUX21X1 U1310 ( .IN1(\regfile[12][31] ), .IN2(AluOut[31]), .S(n1288), .Q(
        n913) );
  MUX21X1 U1311 ( .IN1(\regfile[13][31] ), .IN2(AluOut[31]), .S(n1289), .Q(
        n912) );
  MUX21X1 U1312 ( .IN1(\regfile[14][31] ), .IN2(AluOut[31]), .S(n1290), .Q(
        n911) );
  MUX21X1 U1313 ( .IN1(\regfile[15][31] ), .IN2(AluOut[31]), .S(n1291), .Q(
        n910) );
  AO221X1 U1314 ( .IN1(n1268), .IN2(AluOut[30]), .IN3(N253), .IN4(n1269), 
        .IN5(n1292), .Q(n909) );
  AO21X1 U1315 ( .IN1(n1009), .IN2(IFID_A[30]), .IN3(n1293), .Q(n1292) );
  MUX21X1 U1316 ( .IN1(n1294), .IN2(n1295), .S(IFID_B[30]), .Q(n1293) );
  AO21X1 U1317 ( .IN1(n1274), .IN2(IFID_A[30]), .IN3(n1010), .Q(n1295) );
  NOR2X0 U1318 ( .IN1(n1275), .IN2(IFID_A[30]), .QN(n1294) );
  MUX21X1 U1319 ( .IN1(\regfile[0][30] ), .IN2(AluOut[30]), .S(n1276), .Q(n908) );
  MUX21X1 U1320 ( .IN1(\regfile[1][30] ), .IN2(AluOut[30]), .S(n1277), .Q(n907) );
  MUX21X1 U1321 ( .IN1(\regfile[2][30] ), .IN2(AluOut[30]), .S(n1278), .Q(n906) );
  MUX21X1 U1322 ( .IN1(\regfile[3][30] ), .IN2(AluOut[30]), .S(n1279), .Q(n905) );
  MUX21X1 U1323 ( .IN1(\regfile[4][30] ), .IN2(AluOut[30]), .S(n1280), .Q(n904) );
  MUX21X1 U1324 ( .IN1(\regfile[5][30] ), .IN2(AluOut[30]), .S(n1281), .Q(n903) );
  MUX21X1 U1325 ( .IN1(\regfile[6][30] ), .IN2(AluOut[30]), .S(n1282), .Q(n902) );
  MUX21X1 U1326 ( .IN1(\regfile[7][30] ), .IN2(AluOut[30]), .S(n1283), .Q(n901) );
  MUX21X1 U1327 ( .IN1(\regfile[8][30] ), .IN2(AluOut[30]), .S(n1284), .Q(n900) );
  MUX21X1 U1328 ( .IN1(\regfile[9][30] ), .IN2(AluOut[30]), .S(n1285), .Q(n899) );
  MUX21X1 U1329 ( .IN1(\regfile[10][30] ), .IN2(AluOut[30]), .S(n1286), .Q(
        n898) );
  MUX21X1 U1330 ( .IN1(\regfile[11][30] ), .IN2(AluOut[30]), .S(n1287), .Q(
        n897) );
  MUX21X1 U1331 ( .IN1(\regfile[12][30] ), .IN2(AluOut[30]), .S(n1288), .Q(
        n896) );
  MUX21X1 U1332 ( .IN1(\regfile[13][30] ), .IN2(AluOut[30]), .S(n1289), .Q(
        n895) );
  MUX21X1 U1333 ( .IN1(\regfile[14][30] ), .IN2(AluOut[30]), .S(n1290), .Q(
        n894) );
  MUX21X1 U1334 ( .IN1(\regfile[15][30] ), .IN2(AluOut[30]), .S(n1291), .Q(
        n893) );
  AO221X1 U1335 ( .IN1(n1268), .IN2(AluOut[29]), .IN3(N252), .IN4(n1269), 
        .IN5(n1296), .Q(n892) );
  AO21X1 U1336 ( .IN1(n1008), .IN2(IFID_A[29]), .IN3(n1297), .Q(n1296) );
  MUX21X1 U1337 ( .IN1(n1298), .IN2(n1299), .S(IFID_B[29]), .Q(n1297) );
  AO21X1 U1338 ( .IN1(n1274), .IN2(IFID_A[29]), .IN3(n1009), .Q(n1299) );
  NOR2X0 U1339 ( .IN1(n1275), .IN2(IFID_A[29]), .QN(n1298) );
  MUX21X1 U1340 ( .IN1(\regfile[0][29] ), .IN2(AluOut[29]), .S(n1276), .Q(n891) );
  MUX21X1 U1341 ( .IN1(\regfile[1][29] ), .IN2(AluOut[29]), .S(n1277), .Q(n890) );
  MUX21X1 U1342 ( .IN1(\regfile[2][29] ), .IN2(AluOut[29]), .S(n1278), .Q(n889) );
  MUX21X1 U1343 ( .IN1(\regfile[3][29] ), .IN2(AluOut[29]), .S(n1279), .Q(n888) );
  MUX21X1 U1344 ( .IN1(\regfile[4][29] ), .IN2(AluOut[29]), .S(n1280), .Q(n887) );
  MUX21X1 U1345 ( .IN1(\regfile[5][29] ), .IN2(AluOut[29]), .S(n1281), .Q(n886) );
  MUX21X1 U1346 ( .IN1(\regfile[6][29] ), .IN2(AluOut[29]), .S(n1282), .Q(n885) );
  MUX21X1 U1347 ( .IN1(\regfile[7][29] ), .IN2(AluOut[29]), .S(n1283), .Q(n884) );
  MUX21X1 U1348 ( .IN1(\regfile[8][29] ), .IN2(AluOut[29]), .S(n1284), .Q(n883) );
  MUX21X1 U1349 ( .IN1(\regfile[9][29] ), .IN2(AluOut[29]), .S(n1285), .Q(n882) );
  MUX21X1 U1350 ( .IN1(\regfile[10][29] ), .IN2(AluOut[29]), .S(n1286), .Q(
        n881) );
  MUX21X1 U1351 ( .IN1(\regfile[11][29] ), .IN2(AluOut[29]), .S(n1287), .Q(
        n880) );
  MUX21X1 U1352 ( .IN1(\regfile[12][29] ), .IN2(AluOut[29]), .S(n1288), .Q(
        n879) );
  MUX21X1 U1353 ( .IN1(\regfile[13][29] ), .IN2(AluOut[29]), .S(n1289), .Q(
        n878) );
  MUX21X1 U1354 ( .IN1(\regfile[14][29] ), .IN2(AluOut[29]), .S(n1290), .Q(
        n877) );
  MUX21X1 U1355 ( .IN1(\regfile[15][29] ), .IN2(AluOut[29]), .S(n1291), .Q(
        n876) );
  AO221X1 U1356 ( .IN1(n1268), .IN2(AluOut[28]), .IN3(N251), .IN4(n1269), 
        .IN5(n1300), .Q(n875) );
  AO21X1 U1357 ( .IN1(n1011), .IN2(IFID_A[28]), .IN3(n1301), .Q(n1300) );
  MUX21X1 U1358 ( .IN1(n1302), .IN2(n1303), .S(IFID_B[28]), .Q(n1301) );
  AO21X1 U1359 ( .IN1(n1274), .IN2(IFID_A[28]), .IN3(n1008), .Q(n1303) );
  NOR2X0 U1360 ( .IN1(n1275), .IN2(IFID_A[28]), .QN(n1302) );
  MUX21X1 U1361 ( .IN1(\regfile[0][28] ), .IN2(AluOut[28]), .S(n1276), .Q(n874) );
  MUX21X1 U1362 ( .IN1(\regfile[1][28] ), .IN2(AluOut[28]), .S(n1277), .Q(n873) );
  MUX21X1 U1363 ( .IN1(\regfile[2][28] ), .IN2(AluOut[28]), .S(n1278), .Q(n872) );
  MUX21X1 U1364 ( .IN1(\regfile[3][28] ), .IN2(AluOut[28]), .S(n1279), .Q(n871) );
  MUX21X1 U1365 ( .IN1(\regfile[4][28] ), .IN2(AluOut[28]), .S(n1280), .Q(n870) );
  MUX21X1 U1366 ( .IN1(\regfile[5][28] ), .IN2(AluOut[28]), .S(n1281), .Q(n869) );
  MUX21X1 U1367 ( .IN1(\regfile[6][28] ), .IN2(AluOut[28]), .S(n1282), .Q(n868) );
  MUX21X1 U1368 ( .IN1(\regfile[7][28] ), .IN2(AluOut[28]), .S(n1283), .Q(n867) );
  MUX21X1 U1369 ( .IN1(\regfile[8][28] ), .IN2(AluOut[28]), .S(n1284), .Q(n866) );
  MUX21X1 U1370 ( .IN1(\regfile[9][28] ), .IN2(AluOut[28]), .S(n1285), .Q(n865) );
  MUX21X1 U1371 ( .IN1(\regfile[10][28] ), .IN2(AluOut[28]), .S(n1286), .Q(
        n864) );
  MUX21X1 U1372 ( .IN1(\regfile[11][28] ), .IN2(AluOut[28]), .S(n1287), .Q(
        n863) );
  MUX21X1 U1373 ( .IN1(\regfile[12][28] ), .IN2(AluOut[28]), .S(n1288), .Q(
        n862) );
  MUX21X1 U1374 ( .IN1(\regfile[13][28] ), .IN2(AluOut[28]), .S(n1289), .Q(
        n861) );
  MUX21X1 U1375 ( .IN1(\regfile[14][28] ), .IN2(AluOut[28]), .S(n1290), .Q(
        n860) );
  MUX21X1 U1376 ( .IN1(\regfile[15][28] ), .IN2(AluOut[28]), .S(n1291), .Q(
        n859) );
  AO221X1 U1377 ( .IN1(n1268), .IN2(AluOut[27]), .IN3(N250), .IN4(n1269), 
        .IN5(n1304), .Q(n858) );
  AO21X1 U1378 ( .IN1(n1010), .IN2(IFID_A[27]), .IN3(n1305), .Q(n1304) );
  MUX21X1 U1379 ( .IN1(n1306), .IN2(n1307), .S(IFID_B[27]), .Q(n1305) );
  AO21X1 U1380 ( .IN1(n1274), .IN2(IFID_A[27]), .IN3(n1011), .Q(n1307) );
  NOR2X0 U1381 ( .IN1(n1275), .IN2(IFID_A[27]), .QN(n1306) );
  MUX21X1 U1382 ( .IN1(\regfile[0][27] ), .IN2(AluOut[27]), .S(n1276), .Q(n857) );
  MUX21X1 U1383 ( .IN1(\regfile[1][27] ), .IN2(AluOut[27]), .S(n1277), .Q(n856) );
  MUX21X1 U1384 ( .IN1(\regfile[2][27] ), .IN2(AluOut[27]), .S(n1278), .Q(n855) );
  MUX21X1 U1385 ( .IN1(\regfile[3][27] ), .IN2(AluOut[27]), .S(n1279), .Q(n854) );
  MUX21X1 U1386 ( .IN1(\regfile[4][27] ), .IN2(AluOut[27]), .S(n1280), .Q(n853) );
  MUX21X1 U1387 ( .IN1(\regfile[5][27] ), .IN2(AluOut[27]), .S(n1281), .Q(n852) );
  MUX21X1 U1388 ( .IN1(\regfile[6][27] ), .IN2(AluOut[27]), .S(n1282), .Q(n851) );
  MUX21X1 U1389 ( .IN1(\regfile[7][27] ), .IN2(AluOut[27]), .S(n1283), .Q(n850) );
  MUX21X1 U1390 ( .IN1(\regfile[8][27] ), .IN2(AluOut[27]), .S(n1284), .Q(n849) );
  MUX21X1 U1391 ( .IN1(\regfile[9][27] ), .IN2(AluOut[27]), .S(n1285), .Q(n848) );
  MUX21X1 U1392 ( .IN1(\regfile[10][27] ), .IN2(AluOut[27]), .S(n1286), .Q(
        n847) );
  MUX21X1 U1393 ( .IN1(\regfile[11][27] ), .IN2(AluOut[27]), .S(n1287), .Q(
        n846) );
  MUX21X1 U1394 ( .IN1(\regfile[12][27] ), .IN2(AluOut[27]), .S(n1288), .Q(
        n845) );
  MUX21X1 U1395 ( .IN1(\regfile[13][27] ), .IN2(AluOut[27]), .S(n1289), .Q(
        n844) );
  MUX21X1 U1396 ( .IN1(\regfile[14][27] ), .IN2(AluOut[27]), .S(n1290), .Q(
        n843) );
  MUX21X1 U1397 ( .IN1(\regfile[15][27] ), .IN2(AluOut[27]), .S(n1291), .Q(
        n842) );
  AO221X1 U1398 ( .IN1(n1268), .IN2(AluOut[26]), .IN3(N249), .IN4(n1269), 
        .IN5(n1308), .Q(n841) );
  AO21X1 U1399 ( .IN1(n1009), .IN2(IFID_A[26]), .IN3(n1309), .Q(n1308) );
  MUX21X1 U1400 ( .IN1(n1310), .IN2(n1311), .S(IFID_B[26]), .Q(n1309) );
  AO21X1 U1401 ( .IN1(n1274), .IN2(IFID_A[26]), .IN3(n1010), .Q(n1311) );
  NOR2X0 U1402 ( .IN1(n1275), .IN2(IFID_A[26]), .QN(n1310) );
  MUX21X1 U1403 ( .IN1(\regfile[0][26] ), .IN2(AluOut[26]), .S(n1276), .Q(n840) );
  MUX21X1 U1404 ( .IN1(\regfile[1][26] ), .IN2(AluOut[26]), .S(n1277), .Q(n839) );
  MUX21X1 U1405 ( .IN1(\regfile[2][26] ), .IN2(AluOut[26]), .S(n1278), .Q(n838) );
  MUX21X1 U1406 ( .IN1(\regfile[3][26] ), .IN2(AluOut[26]), .S(n1279), .Q(n837) );
  MUX21X1 U1407 ( .IN1(\regfile[4][26] ), .IN2(AluOut[26]), .S(n1280), .Q(n836) );
  MUX21X1 U1408 ( .IN1(\regfile[5][26] ), .IN2(AluOut[26]), .S(n1281), .Q(n835) );
  MUX21X1 U1409 ( .IN1(\regfile[6][26] ), .IN2(AluOut[26]), .S(n1282), .Q(n834) );
  MUX21X1 U1410 ( .IN1(\regfile[7][26] ), .IN2(AluOut[26]), .S(n1283), .Q(n833) );
  MUX21X1 U1411 ( .IN1(\regfile[8][26] ), .IN2(AluOut[26]), .S(n1284), .Q(n832) );
  MUX21X1 U1412 ( .IN1(\regfile[9][26] ), .IN2(AluOut[26]), .S(n1285), .Q(n831) );
  MUX21X1 U1413 ( .IN1(\regfile[10][26] ), .IN2(AluOut[26]), .S(n1286), .Q(
        n830) );
  MUX21X1 U1414 ( .IN1(\regfile[11][26] ), .IN2(AluOut[26]), .S(n1287), .Q(
        n829) );
  MUX21X1 U1415 ( .IN1(\regfile[12][26] ), .IN2(AluOut[26]), .S(n1288), .Q(
        n828) );
  MUX21X1 U1416 ( .IN1(\regfile[13][26] ), .IN2(AluOut[26]), .S(n1289), .Q(
        n827) );
  MUX21X1 U1417 ( .IN1(\regfile[14][26] ), .IN2(AluOut[26]), .S(n1290), .Q(
        n826) );
  MUX21X1 U1418 ( .IN1(\regfile[15][26] ), .IN2(AluOut[26]), .S(n1291), .Q(
        n825) );
  AO221X1 U1419 ( .IN1(n1268), .IN2(AluOut[25]), .IN3(N248), .IN4(n1269), 
        .IN5(n1312), .Q(n824) );
  AO21X1 U1420 ( .IN1(n1008), .IN2(IFID_A[25]), .IN3(n1313), .Q(n1312) );
  MUX21X1 U1421 ( .IN1(n1314), .IN2(n1315), .S(IFID_B[25]), .Q(n1313) );
  AO21X1 U1422 ( .IN1(n1274), .IN2(IFID_A[25]), .IN3(n1009), .Q(n1315) );
  NOR2X0 U1423 ( .IN1(n1275), .IN2(IFID_A[25]), .QN(n1314) );
  MUX21X1 U1424 ( .IN1(\regfile[0][25] ), .IN2(AluOut[25]), .S(n1276), .Q(n823) );
  MUX21X1 U1425 ( .IN1(\regfile[1][25] ), .IN2(AluOut[25]), .S(n1277), .Q(n822) );
  MUX21X1 U1426 ( .IN1(\regfile[2][25] ), .IN2(AluOut[25]), .S(n1278), .Q(n821) );
  MUX21X1 U1427 ( .IN1(\regfile[3][25] ), .IN2(AluOut[25]), .S(n1279), .Q(n820) );
  MUX21X1 U1428 ( .IN1(\regfile[4][25] ), .IN2(AluOut[25]), .S(n1280), .Q(n819) );
  MUX21X1 U1429 ( .IN1(\regfile[5][25] ), .IN2(AluOut[25]), .S(n1281), .Q(n818) );
  MUX21X1 U1430 ( .IN1(\regfile[6][25] ), .IN2(AluOut[25]), .S(n1282), .Q(n817) );
  MUX21X1 U1431 ( .IN1(\regfile[7][25] ), .IN2(AluOut[25]), .S(n1283), .Q(n816) );
  MUX21X1 U1432 ( .IN1(\regfile[8][25] ), .IN2(AluOut[25]), .S(n1284), .Q(n815) );
  MUX21X1 U1433 ( .IN1(\regfile[9][25] ), .IN2(AluOut[25]), .S(n1285), .Q(n814) );
  MUX21X1 U1434 ( .IN1(\regfile[10][25] ), .IN2(AluOut[25]), .S(n1286), .Q(
        n813) );
  MUX21X1 U1435 ( .IN1(\regfile[11][25] ), .IN2(AluOut[25]), .S(n1287), .Q(
        n812) );
  MUX21X1 U1436 ( .IN1(\regfile[12][25] ), .IN2(AluOut[25]), .S(n1288), .Q(
        n811) );
  MUX21X1 U1437 ( .IN1(\regfile[13][25] ), .IN2(AluOut[25]), .S(n1289), .Q(
        n810) );
  MUX21X1 U1438 ( .IN1(\regfile[14][25] ), .IN2(AluOut[25]), .S(n1290), .Q(
        n809) );
  MUX21X1 U1439 ( .IN1(\regfile[15][25] ), .IN2(AluOut[25]), .S(n1291), .Q(
        n808) );
  AO221X1 U1440 ( .IN1(n1268), .IN2(AluOut[24]), .IN3(N247), .IN4(n1269), 
        .IN5(n1316), .Q(n807) );
  AO21X1 U1441 ( .IN1(n1011), .IN2(IFID_A[24]), .IN3(n1317), .Q(n1316) );
  MUX21X1 U1442 ( .IN1(n1318), .IN2(n1319), .S(IFID_B[24]), .Q(n1317) );
  AO21X1 U1443 ( .IN1(n1274), .IN2(IFID_A[24]), .IN3(n1008), .Q(n1319) );
  NOR2X0 U1444 ( .IN1(n1275), .IN2(IFID_A[24]), .QN(n1318) );
  MUX21X1 U1445 ( .IN1(\regfile[0][24] ), .IN2(AluOut[24]), .S(n1276), .Q(n806) );
  MUX21X1 U1446 ( .IN1(\regfile[1][24] ), .IN2(AluOut[24]), .S(n1277), .Q(n805) );
  MUX21X1 U1447 ( .IN1(\regfile[2][24] ), .IN2(AluOut[24]), .S(n1278), .Q(n804) );
  MUX21X1 U1448 ( .IN1(\regfile[3][24] ), .IN2(AluOut[24]), .S(n1279), .Q(n803) );
  MUX21X1 U1449 ( .IN1(\regfile[4][24] ), .IN2(AluOut[24]), .S(n1280), .Q(n802) );
  MUX21X1 U1450 ( .IN1(\regfile[5][24] ), .IN2(AluOut[24]), .S(n1281), .Q(n801) );
  MUX21X1 U1451 ( .IN1(\regfile[6][24] ), .IN2(AluOut[24]), .S(n1282), .Q(n800) );
  MUX21X1 U1452 ( .IN1(\regfile[7][24] ), .IN2(AluOut[24]), .S(n1283), .Q(n799) );
  MUX21X1 U1453 ( .IN1(\regfile[8][24] ), .IN2(AluOut[24]), .S(n1284), .Q(n798) );
  MUX21X1 U1454 ( .IN1(\regfile[9][24] ), .IN2(AluOut[24]), .S(n1285), .Q(n797) );
  MUX21X1 U1455 ( .IN1(\regfile[10][24] ), .IN2(AluOut[24]), .S(n1286), .Q(
        n796) );
  MUX21X1 U1456 ( .IN1(\regfile[11][24] ), .IN2(AluOut[24]), .S(n1287), .Q(
        n795) );
  MUX21X1 U1457 ( .IN1(\regfile[12][24] ), .IN2(AluOut[24]), .S(n1288), .Q(
        n794) );
  MUX21X1 U1458 ( .IN1(\regfile[13][24] ), .IN2(AluOut[24]), .S(n1289), .Q(
        n793) );
  MUX21X1 U1459 ( .IN1(\regfile[14][24] ), .IN2(AluOut[24]), .S(n1290), .Q(
        n792) );
  MUX21X1 U1460 ( .IN1(\regfile[15][24] ), .IN2(AluOut[24]), .S(n1291), .Q(
        n791) );
  AO221X1 U1461 ( .IN1(n1268), .IN2(AluOut[23]), .IN3(N246), .IN4(n1269), 
        .IN5(n1320), .Q(n790) );
  AO21X1 U1462 ( .IN1(n1010), .IN2(IFID_A[23]), .IN3(n1321), .Q(n1320) );
  MUX21X1 U1463 ( .IN1(n1322), .IN2(n1323), .S(IFID_B[23]), .Q(n1321) );
  AO21X1 U1464 ( .IN1(n1274), .IN2(IFID_A[23]), .IN3(n1011), .Q(n1323) );
  NOR2X0 U1465 ( .IN1(n1275), .IN2(IFID_A[23]), .QN(n1322) );
  MUX21X1 U1466 ( .IN1(\regfile[0][23] ), .IN2(AluOut[23]), .S(n1276), .Q(n789) );
  MUX21X1 U1467 ( .IN1(\regfile[1][23] ), .IN2(AluOut[23]), .S(n1277), .Q(n788) );
  MUX21X1 U1468 ( .IN1(\regfile[2][23] ), .IN2(AluOut[23]), .S(n1278), .Q(n787) );
  MUX21X1 U1469 ( .IN1(\regfile[3][23] ), .IN2(AluOut[23]), .S(n1279), .Q(n786) );
  MUX21X1 U1470 ( .IN1(\regfile[4][23] ), .IN2(AluOut[23]), .S(n1280), .Q(n785) );
  MUX21X1 U1471 ( .IN1(\regfile[5][23] ), .IN2(AluOut[23]), .S(n1281), .Q(n784) );
  MUX21X1 U1472 ( .IN1(\regfile[6][23] ), .IN2(AluOut[23]), .S(n1282), .Q(n783) );
  MUX21X1 U1473 ( .IN1(\regfile[7][23] ), .IN2(AluOut[23]), .S(n1283), .Q(n782) );
  MUX21X1 U1474 ( .IN1(\regfile[8][23] ), .IN2(AluOut[23]), .S(n1284), .Q(n781) );
  MUX21X1 U1475 ( .IN1(\regfile[9][23] ), .IN2(AluOut[23]), .S(n1285), .Q(n780) );
  MUX21X1 U1476 ( .IN1(\regfile[10][23] ), .IN2(AluOut[23]), .S(n1286), .Q(
        n779) );
  MUX21X1 U1477 ( .IN1(\regfile[11][23] ), .IN2(AluOut[23]), .S(n1287), .Q(
        n778) );
  MUX21X1 U1478 ( .IN1(\regfile[12][23] ), .IN2(AluOut[23]), .S(n1288), .Q(
        n777) );
  MUX21X1 U1479 ( .IN1(\regfile[13][23] ), .IN2(AluOut[23]), .S(n1289), .Q(
        n776) );
  MUX21X1 U1480 ( .IN1(\regfile[14][23] ), .IN2(AluOut[23]), .S(n1290), .Q(
        n775) );
  MUX21X1 U1481 ( .IN1(\regfile[15][23] ), .IN2(AluOut[23]), .S(n1291), .Q(
        n774) );
  AO221X1 U1482 ( .IN1(n1268), .IN2(AluOut[22]), .IN3(N245), .IN4(n1269), 
        .IN5(n1324), .Q(n773) );
  AO21X1 U1483 ( .IN1(n1009), .IN2(IFID_A[22]), .IN3(n1325), .Q(n1324) );
  MUX21X1 U1484 ( .IN1(n1326), .IN2(n1327), .S(IFID_B[22]), .Q(n1325) );
  AO21X1 U1485 ( .IN1(n1274), .IN2(IFID_A[22]), .IN3(n1010), .Q(n1327) );
  NOR2X0 U1486 ( .IN1(n1275), .IN2(IFID_A[22]), .QN(n1326) );
  MUX21X1 U1487 ( .IN1(\regfile[0][22] ), .IN2(AluOut[22]), .S(n1276), .Q(n772) );
  MUX21X1 U1488 ( .IN1(\regfile[1][22] ), .IN2(AluOut[22]), .S(n1277), .Q(n771) );
  MUX21X1 U1489 ( .IN1(\regfile[2][22] ), .IN2(AluOut[22]), .S(n1278), .Q(n770) );
  MUX21X1 U1490 ( .IN1(\regfile[3][22] ), .IN2(AluOut[22]), .S(n1279), .Q(n769) );
  MUX21X1 U1491 ( .IN1(\regfile[4][22] ), .IN2(AluOut[22]), .S(n1280), .Q(n768) );
  MUX21X1 U1492 ( .IN1(\regfile[5][22] ), .IN2(AluOut[22]), .S(n1281), .Q(n767) );
  MUX21X1 U1493 ( .IN1(\regfile[6][22] ), .IN2(AluOut[22]), .S(n1282), .Q(n766) );
  MUX21X1 U1494 ( .IN1(\regfile[7][22] ), .IN2(AluOut[22]), .S(n1283), .Q(n765) );
  MUX21X1 U1495 ( .IN1(\regfile[8][22] ), .IN2(AluOut[22]), .S(n1284), .Q(n764) );
  MUX21X1 U1496 ( .IN1(\regfile[9][22] ), .IN2(AluOut[22]), .S(n1285), .Q(n763) );
  MUX21X1 U1497 ( .IN1(\regfile[10][22] ), .IN2(AluOut[22]), .S(n1286), .Q(
        n762) );
  MUX21X1 U1498 ( .IN1(\regfile[11][22] ), .IN2(AluOut[22]), .S(n1287), .Q(
        n761) );
  MUX21X1 U1499 ( .IN1(\regfile[12][22] ), .IN2(AluOut[22]), .S(n1288), .Q(
        n760) );
  MUX21X1 U1500 ( .IN1(\regfile[13][22] ), .IN2(AluOut[22]), .S(n1289), .Q(
        n759) );
  MUX21X1 U1501 ( .IN1(\regfile[14][22] ), .IN2(AluOut[22]), .S(n1290), .Q(
        n758) );
  MUX21X1 U1502 ( .IN1(\regfile[15][22] ), .IN2(AluOut[22]), .S(n1291), .Q(
        n757) );
  AO221X1 U1503 ( .IN1(n1268), .IN2(AluOut[21]), .IN3(N244), .IN4(n1269), 
        .IN5(n1328), .Q(n756) );
  AO21X1 U1504 ( .IN1(n1008), .IN2(IFID_A[21]), .IN3(n1329), .Q(n1328) );
  MUX21X1 U1505 ( .IN1(n1330), .IN2(n1331), .S(IFID_B[21]), .Q(n1329) );
  AO21X1 U1506 ( .IN1(n1274), .IN2(IFID_A[21]), .IN3(n1009), .Q(n1331) );
  NOR2X0 U1507 ( .IN1(n1275), .IN2(IFID_A[21]), .QN(n1330) );
  MUX21X1 U1508 ( .IN1(\regfile[0][21] ), .IN2(AluOut[21]), .S(n1276), .Q(n755) );
  MUX21X1 U1509 ( .IN1(\regfile[1][21] ), .IN2(AluOut[21]), .S(n1277), .Q(n754) );
  MUX21X1 U1510 ( .IN1(\regfile[2][21] ), .IN2(AluOut[21]), .S(n1278), .Q(n753) );
  MUX21X1 U1511 ( .IN1(\regfile[3][21] ), .IN2(AluOut[21]), .S(n1279), .Q(n752) );
  MUX21X1 U1512 ( .IN1(\regfile[4][21] ), .IN2(AluOut[21]), .S(n1280), .Q(n751) );
  MUX21X1 U1513 ( .IN1(\regfile[5][21] ), .IN2(AluOut[21]), .S(n1281), .Q(n750) );
  MUX21X1 U1514 ( .IN1(\regfile[6][21] ), .IN2(AluOut[21]), .S(n1282), .Q(n749) );
  MUX21X1 U1515 ( .IN1(\regfile[7][21] ), .IN2(AluOut[21]), .S(n1283), .Q(n748) );
  MUX21X1 U1516 ( .IN1(\regfile[8][21] ), .IN2(AluOut[21]), .S(n1284), .Q(n747) );
  MUX21X1 U1517 ( .IN1(\regfile[9][21] ), .IN2(AluOut[21]), .S(n1285), .Q(n746) );
  MUX21X1 U1518 ( .IN1(\regfile[10][21] ), .IN2(AluOut[21]), .S(n1286), .Q(
        n745) );
  MUX21X1 U1519 ( .IN1(\regfile[11][21] ), .IN2(AluOut[21]), .S(n1287), .Q(
        n744) );
  MUX21X1 U1520 ( .IN1(\regfile[12][21] ), .IN2(AluOut[21]), .S(n1288), .Q(
        n743) );
  MUX21X1 U1521 ( .IN1(\regfile[13][21] ), .IN2(AluOut[21]), .S(n1289), .Q(
        n742) );
  MUX21X1 U1522 ( .IN1(\regfile[14][21] ), .IN2(AluOut[21]), .S(n1290), .Q(
        n741) );
  MUX21X1 U1523 ( .IN1(\regfile[15][21] ), .IN2(AluOut[21]), .S(n1291), .Q(
        n740) );
  AO221X1 U1524 ( .IN1(n1268), .IN2(AluOut[20]), .IN3(N243), .IN4(n1269), 
        .IN5(n1332), .Q(n739) );
  AO21X1 U1525 ( .IN1(n1011), .IN2(IFID_A[20]), .IN3(n1333), .Q(n1332) );
  MUX21X1 U1526 ( .IN1(n1334), .IN2(n1335), .S(IFID_B[20]), .Q(n1333) );
  AO21X1 U1527 ( .IN1(n1274), .IN2(IFID_A[20]), .IN3(n1008), .Q(n1335) );
  NOR2X0 U1528 ( .IN1(n1275), .IN2(IFID_A[20]), .QN(n1334) );
  MUX21X1 U1529 ( .IN1(\regfile[0][20] ), .IN2(AluOut[20]), .S(n1276), .Q(n738) );
  MUX21X1 U1530 ( .IN1(\regfile[1][20] ), .IN2(AluOut[20]), .S(n1277), .Q(n737) );
  MUX21X1 U1531 ( .IN1(\regfile[2][20] ), .IN2(AluOut[20]), .S(n1278), .Q(n736) );
  MUX21X1 U1532 ( .IN1(\regfile[3][20] ), .IN2(AluOut[20]), .S(n1279), .Q(n735) );
  MUX21X1 U1533 ( .IN1(\regfile[4][20] ), .IN2(AluOut[20]), .S(n1280), .Q(n734) );
  MUX21X1 U1534 ( .IN1(\regfile[5][20] ), .IN2(AluOut[20]), .S(n1281), .Q(n733) );
  MUX21X1 U1535 ( .IN1(\regfile[6][20] ), .IN2(AluOut[20]), .S(n1282), .Q(n732) );
  MUX21X1 U1536 ( .IN1(\regfile[7][20] ), .IN2(AluOut[20]), .S(n1283), .Q(n731) );
  MUX21X1 U1537 ( .IN1(\regfile[8][20] ), .IN2(AluOut[20]), .S(n1284), .Q(n730) );
  MUX21X1 U1538 ( .IN1(\regfile[9][20] ), .IN2(AluOut[20]), .S(n1285), .Q(n729) );
  MUX21X1 U1539 ( .IN1(\regfile[10][20] ), .IN2(AluOut[20]), .S(n1286), .Q(
        n728) );
  MUX21X1 U1540 ( .IN1(\regfile[11][20] ), .IN2(AluOut[20]), .S(n1287), .Q(
        n727) );
  MUX21X1 U1541 ( .IN1(\regfile[12][20] ), .IN2(AluOut[20]), .S(n1288), .Q(
        n726) );
  MUX21X1 U1542 ( .IN1(\regfile[13][20] ), .IN2(AluOut[20]), .S(n1289), .Q(
        n725) );
  MUX21X1 U1543 ( .IN1(\regfile[14][20] ), .IN2(AluOut[20]), .S(n1290), .Q(
        n724) );
  MUX21X1 U1544 ( .IN1(\regfile[15][20] ), .IN2(AluOut[20]), .S(n1291), .Q(
        n723) );
  AO221X1 U1545 ( .IN1(n1268), .IN2(AluOut[19]), .IN3(N242), .IN4(n1269), 
        .IN5(n1336), .Q(n722) );
  AO21X1 U1546 ( .IN1(n1010), .IN2(IFID_A[19]), .IN3(n1337), .Q(n1336) );
  MUX21X1 U1547 ( .IN1(n1338), .IN2(n1339), .S(IFID_B[19]), .Q(n1337) );
  AO21X1 U1548 ( .IN1(n1274), .IN2(IFID_A[19]), .IN3(n1011), .Q(n1339) );
  NOR2X0 U1549 ( .IN1(n1275), .IN2(IFID_A[19]), .QN(n1338) );
  MUX21X1 U1550 ( .IN1(\regfile[0][19] ), .IN2(AluOut[19]), .S(n1276), .Q(n721) );
  MUX21X1 U1551 ( .IN1(\regfile[1][19] ), .IN2(AluOut[19]), .S(n1277), .Q(n720) );
  MUX21X1 U1552 ( .IN1(\regfile[2][19] ), .IN2(AluOut[19]), .S(n1278), .Q(n719) );
  MUX21X1 U1553 ( .IN1(\regfile[3][19] ), .IN2(AluOut[19]), .S(n1279), .Q(n718) );
  MUX21X1 U1554 ( .IN1(\regfile[4][19] ), .IN2(AluOut[19]), .S(n1280), .Q(n717) );
  MUX21X1 U1555 ( .IN1(\regfile[5][19] ), .IN2(AluOut[19]), .S(n1281), .Q(n716) );
  MUX21X1 U1556 ( .IN1(\regfile[6][19] ), .IN2(AluOut[19]), .S(n1282), .Q(n715) );
  MUX21X1 U1557 ( .IN1(\regfile[7][19] ), .IN2(AluOut[19]), .S(n1283), .Q(n714) );
  MUX21X1 U1558 ( .IN1(\regfile[8][19] ), .IN2(AluOut[19]), .S(n1284), .Q(n713) );
  MUX21X1 U1559 ( .IN1(\regfile[9][19] ), .IN2(AluOut[19]), .S(n1285), .Q(n712) );
  MUX21X1 U1560 ( .IN1(\regfile[10][19] ), .IN2(AluOut[19]), .S(n1286), .Q(
        n711) );
  MUX21X1 U1561 ( .IN1(\regfile[11][19] ), .IN2(AluOut[19]), .S(n1287), .Q(
        n710) );
  MUX21X1 U1562 ( .IN1(\regfile[12][19] ), .IN2(AluOut[19]), .S(n1288), .Q(
        n709) );
  MUX21X1 U1563 ( .IN1(\regfile[13][19] ), .IN2(AluOut[19]), .S(n1289), .Q(
        n708) );
  MUX21X1 U1564 ( .IN1(\regfile[14][19] ), .IN2(AluOut[19]), .S(n1290), .Q(
        n707) );
  MUX21X1 U1565 ( .IN1(\regfile[15][19] ), .IN2(AluOut[19]), .S(n1291), .Q(
        n706) );
  AO221X1 U1566 ( .IN1(n1268), .IN2(AluOut[18]), .IN3(N241), .IN4(n1269), 
        .IN5(n1340), .Q(n705) );
  AO21X1 U1567 ( .IN1(n1009), .IN2(IFID_A[18]), .IN3(n1341), .Q(n1340) );
  MUX21X1 U1568 ( .IN1(n1342), .IN2(n1343), .S(IFID_B[18]), .Q(n1341) );
  AO21X1 U1569 ( .IN1(n1274), .IN2(IFID_A[18]), .IN3(n1010), .Q(n1343) );
  NOR2X0 U1570 ( .IN1(n1275), .IN2(IFID_A[18]), .QN(n1342) );
  MUX21X1 U1571 ( .IN1(\regfile[0][18] ), .IN2(AluOut[18]), .S(n1276), .Q(n704) );
  MUX21X1 U1572 ( .IN1(\regfile[1][18] ), .IN2(AluOut[18]), .S(n1277), .Q(n703) );
  MUX21X1 U1573 ( .IN1(\regfile[2][18] ), .IN2(AluOut[18]), .S(n1278), .Q(n702) );
  MUX21X1 U1574 ( .IN1(\regfile[3][18] ), .IN2(AluOut[18]), .S(n1279), .Q(n701) );
  MUX21X1 U1575 ( .IN1(\regfile[4][18] ), .IN2(AluOut[18]), .S(n1280), .Q(n700) );
  MUX21X1 U1576 ( .IN1(\regfile[5][18] ), .IN2(AluOut[18]), .S(n1281), .Q(n699) );
  MUX21X1 U1577 ( .IN1(\regfile[6][18] ), .IN2(AluOut[18]), .S(n1282), .Q(n698) );
  MUX21X1 U1578 ( .IN1(\regfile[7][18] ), .IN2(AluOut[18]), .S(n1283), .Q(n697) );
  MUX21X1 U1579 ( .IN1(\regfile[8][18] ), .IN2(AluOut[18]), .S(n1284), .Q(n696) );
  MUX21X1 U1580 ( .IN1(\regfile[9][18] ), .IN2(AluOut[18]), .S(n1285), .Q(n695) );
  MUX21X1 U1581 ( .IN1(\regfile[10][18] ), .IN2(AluOut[18]), .S(n1286), .Q(
        n694) );
  MUX21X1 U1582 ( .IN1(\regfile[11][18] ), .IN2(AluOut[18]), .S(n1287), .Q(
        n693) );
  MUX21X1 U1583 ( .IN1(\regfile[12][18] ), .IN2(AluOut[18]), .S(n1288), .Q(
        n692) );
  MUX21X1 U1584 ( .IN1(\regfile[13][18] ), .IN2(AluOut[18]), .S(n1289), .Q(
        n691) );
  MUX21X1 U1585 ( .IN1(\regfile[14][18] ), .IN2(AluOut[18]), .S(n1290), .Q(
        n690) );
  MUX21X1 U1586 ( .IN1(\regfile[15][18] ), .IN2(AluOut[18]), .S(n1291), .Q(
        n689) );
  AO221X1 U1587 ( .IN1(n1268), .IN2(AluOut[17]), .IN3(N240), .IN4(n1269), 
        .IN5(n1344), .Q(n688) );
  AO21X1 U1588 ( .IN1(n1008), .IN2(IFID_A[17]), .IN3(n1345), .Q(n1344) );
  MUX21X1 U1589 ( .IN1(n1346), .IN2(n1347), .S(IFID_B[17]), .Q(n1345) );
  AO21X1 U1590 ( .IN1(n1274), .IN2(IFID_A[17]), .IN3(n1009), .Q(n1347) );
  NOR2X0 U1591 ( .IN1(n1275), .IN2(IFID_A[17]), .QN(n1346) );
  MUX21X1 U1592 ( .IN1(\regfile[0][17] ), .IN2(AluOut[17]), .S(n1276), .Q(n687) );
  MUX21X1 U1593 ( .IN1(\regfile[1][17] ), .IN2(AluOut[17]), .S(n1277), .Q(n686) );
  MUX21X1 U1594 ( .IN1(\regfile[2][17] ), .IN2(AluOut[17]), .S(n1278), .Q(n685) );
  MUX21X1 U1595 ( .IN1(\regfile[3][17] ), .IN2(AluOut[17]), .S(n1279), .Q(n684) );
  MUX21X1 U1596 ( .IN1(\regfile[4][17] ), .IN2(AluOut[17]), .S(n1280), .Q(n683) );
  MUX21X1 U1597 ( .IN1(\regfile[5][17] ), .IN2(AluOut[17]), .S(n1281), .Q(n682) );
  MUX21X1 U1598 ( .IN1(\regfile[6][17] ), .IN2(AluOut[17]), .S(n1282), .Q(n681) );
  MUX21X1 U1599 ( .IN1(\regfile[7][17] ), .IN2(AluOut[17]), .S(n1283), .Q(n680) );
  MUX21X1 U1600 ( .IN1(\regfile[8][17] ), .IN2(AluOut[17]), .S(n1284), .Q(n679) );
  MUX21X1 U1601 ( .IN1(\regfile[9][17] ), .IN2(AluOut[17]), .S(n1285), .Q(n678) );
  MUX21X1 U1602 ( .IN1(\regfile[10][17] ), .IN2(AluOut[17]), .S(n1286), .Q(
        n677) );
  MUX21X1 U1603 ( .IN1(\regfile[11][17] ), .IN2(AluOut[17]), .S(n1287), .Q(
        n676) );
  MUX21X1 U1604 ( .IN1(\regfile[12][17] ), .IN2(AluOut[17]), .S(n1288), .Q(
        n675) );
  MUX21X1 U1605 ( .IN1(\regfile[13][17] ), .IN2(AluOut[17]), .S(n1289), .Q(
        n674) );
  MUX21X1 U1606 ( .IN1(\regfile[14][17] ), .IN2(AluOut[17]), .S(n1290), .Q(
        n673) );
  MUX21X1 U1607 ( .IN1(\regfile[15][17] ), .IN2(AluOut[17]), .S(n1291), .Q(
        n672) );
  AO221X1 U1608 ( .IN1(n1268), .IN2(AluOut[16]), .IN3(N239), .IN4(n1269), 
        .IN5(n1348), .Q(n671) );
  AO21X1 U1609 ( .IN1(n1011), .IN2(IFID_A[16]), .IN3(n1349), .Q(n1348) );
  MUX21X1 U1610 ( .IN1(n1350), .IN2(n1351), .S(IFID_B[16]), .Q(n1349) );
  AO21X1 U1611 ( .IN1(n1274), .IN2(IFID_A[16]), .IN3(n1008), .Q(n1351) );
  NOR2X0 U1612 ( .IN1(n1275), .IN2(IFID_A[16]), .QN(n1350) );
  MUX21X1 U1613 ( .IN1(\regfile[0][16] ), .IN2(AluOut[16]), .S(n1276), .Q(n670) );
  MUX21X1 U1614 ( .IN1(\regfile[1][16] ), .IN2(AluOut[16]), .S(n1277), .Q(n669) );
  MUX21X1 U1615 ( .IN1(\regfile[2][16] ), .IN2(AluOut[16]), .S(n1278), .Q(n668) );
  MUX21X1 U1616 ( .IN1(\regfile[3][16] ), .IN2(AluOut[16]), .S(n1279), .Q(n667) );
  MUX21X1 U1617 ( .IN1(\regfile[4][16] ), .IN2(AluOut[16]), .S(n1280), .Q(n666) );
  MUX21X1 U1618 ( .IN1(\regfile[5][16] ), .IN2(AluOut[16]), .S(n1281), .Q(n665) );
  MUX21X1 U1619 ( .IN1(\regfile[6][16] ), .IN2(AluOut[16]), .S(n1282), .Q(n664) );
  MUX21X1 U1620 ( .IN1(\regfile[7][16] ), .IN2(AluOut[16]), .S(n1283), .Q(n663) );
  MUX21X1 U1621 ( .IN1(\regfile[8][16] ), .IN2(AluOut[16]), .S(n1284), .Q(n662) );
  MUX21X1 U1622 ( .IN1(\regfile[9][16] ), .IN2(AluOut[16]), .S(n1285), .Q(n661) );
  MUX21X1 U1623 ( .IN1(\regfile[10][16] ), .IN2(AluOut[16]), .S(n1286), .Q(
        n660) );
  MUX21X1 U1624 ( .IN1(\regfile[11][16] ), .IN2(AluOut[16]), .S(n1287), .Q(
        n659) );
  MUX21X1 U1625 ( .IN1(\regfile[12][16] ), .IN2(AluOut[16]), .S(n1288), .Q(
        n658) );
  MUX21X1 U1626 ( .IN1(\regfile[13][16] ), .IN2(AluOut[16]), .S(n1289), .Q(
        n657) );
  MUX21X1 U1627 ( .IN1(\regfile[14][16] ), .IN2(AluOut[16]), .S(n1290), .Q(
        n656) );
  MUX21X1 U1628 ( .IN1(\regfile[15][16] ), .IN2(AluOut[16]), .S(n1291), .Q(
        n655) );
  AO221X1 U1629 ( .IN1(n1268), .IN2(AluOut[15]), .IN3(N238), .IN4(n1269), 
        .IN5(n1352), .Q(n654) );
  AO21X1 U1630 ( .IN1(n1010), .IN2(IFID_A[15]), .IN3(n1353), .Q(n1352) );
  MUX21X1 U1631 ( .IN1(n1354), .IN2(n1355), .S(IFID_B[15]), .Q(n1353) );
  AO21X1 U1632 ( .IN1(n1274), .IN2(IFID_A[15]), .IN3(n1011), .Q(n1355) );
  NOR2X0 U1633 ( .IN1(n1275), .IN2(IFID_A[15]), .QN(n1354) );
  MUX21X1 U1634 ( .IN1(\regfile[0][15] ), .IN2(AluOut[15]), .S(n1276), .Q(n653) );
  MUX21X1 U1635 ( .IN1(\regfile[1][15] ), .IN2(AluOut[15]), .S(n1277), .Q(n652) );
  MUX21X1 U1636 ( .IN1(\regfile[2][15] ), .IN2(AluOut[15]), .S(n1278), .Q(n651) );
  MUX21X1 U1637 ( .IN1(\regfile[3][15] ), .IN2(AluOut[15]), .S(n1279), .Q(n650) );
  MUX21X1 U1638 ( .IN1(\regfile[4][15] ), .IN2(AluOut[15]), .S(n1280), .Q(n649) );
  MUX21X1 U1639 ( .IN1(\regfile[5][15] ), .IN2(AluOut[15]), .S(n1281), .Q(n648) );
  MUX21X1 U1640 ( .IN1(\regfile[6][15] ), .IN2(AluOut[15]), .S(n1282), .Q(n647) );
  MUX21X1 U1641 ( .IN1(\regfile[7][15] ), .IN2(AluOut[15]), .S(n1283), .Q(n646) );
  MUX21X1 U1642 ( .IN1(\regfile[8][15] ), .IN2(AluOut[15]), .S(n1284), .Q(n645) );
  MUX21X1 U1643 ( .IN1(\regfile[9][15] ), .IN2(AluOut[15]), .S(n1285), .Q(n644) );
  MUX21X1 U1644 ( .IN1(\regfile[10][15] ), .IN2(AluOut[15]), .S(n1286), .Q(
        n643) );
  MUX21X1 U1645 ( .IN1(\regfile[11][15] ), .IN2(AluOut[15]), .S(n1287), .Q(
        n642) );
  MUX21X1 U1646 ( .IN1(\regfile[12][15] ), .IN2(AluOut[15]), .S(n1288), .Q(
        n641) );
  MUX21X1 U1647 ( .IN1(\regfile[13][15] ), .IN2(AluOut[15]), .S(n1289), .Q(
        n640) );
  MUX21X1 U1648 ( .IN1(\regfile[14][15] ), .IN2(AluOut[15]), .S(n1290), .Q(
        n639) );
  MUX21X1 U1649 ( .IN1(\regfile[15][15] ), .IN2(AluOut[15]), .S(n1291), .Q(
        n638) );
  AO221X1 U1650 ( .IN1(n1268), .IN2(AluOut[14]), .IN3(N237), .IN4(n1269), 
        .IN5(n1356), .Q(n637) );
  AO21X1 U1651 ( .IN1(n1009), .IN2(IFID_A[14]), .IN3(n1357), .Q(n1356) );
  MUX21X1 U1652 ( .IN1(n1358), .IN2(n1359), .S(IFID_B[14]), .Q(n1357) );
  AO21X1 U1653 ( .IN1(n1274), .IN2(IFID_A[14]), .IN3(n1010), .Q(n1359) );
  NOR2X0 U1654 ( .IN1(n1275), .IN2(IFID_A[14]), .QN(n1358) );
  MUX21X1 U1655 ( .IN1(\regfile[0][14] ), .IN2(AluOut[14]), .S(n1276), .Q(n636) );
  MUX21X1 U1656 ( .IN1(\regfile[1][14] ), .IN2(AluOut[14]), .S(n1277), .Q(n635) );
  MUX21X1 U1657 ( .IN1(\regfile[2][14] ), .IN2(AluOut[14]), .S(n1278), .Q(n634) );
  MUX21X1 U1658 ( .IN1(\regfile[3][14] ), .IN2(AluOut[14]), .S(n1279), .Q(n633) );
  MUX21X1 U1659 ( .IN1(\regfile[4][14] ), .IN2(AluOut[14]), .S(n1280), .Q(n632) );
  MUX21X1 U1660 ( .IN1(\regfile[5][14] ), .IN2(AluOut[14]), .S(n1281), .Q(n631) );
  MUX21X1 U1661 ( .IN1(\regfile[6][14] ), .IN2(AluOut[14]), .S(n1282), .Q(n630) );
  MUX21X1 U1662 ( .IN1(\regfile[7][14] ), .IN2(AluOut[14]), .S(n1283), .Q(n629) );
  MUX21X1 U1663 ( .IN1(\regfile[8][14] ), .IN2(AluOut[14]), .S(n1284), .Q(n628) );
  MUX21X1 U1664 ( .IN1(\regfile[9][14] ), .IN2(AluOut[14]), .S(n1285), .Q(n627) );
  MUX21X1 U1665 ( .IN1(\regfile[10][14] ), .IN2(AluOut[14]), .S(n1286), .Q(
        n626) );
  MUX21X1 U1666 ( .IN1(\regfile[11][14] ), .IN2(AluOut[14]), .S(n1287), .Q(
        n625) );
  MUX21X1 U1667 ( .IN1(\regfile[12][14] ), .IN2(AluOut[14]), .S(n1288), .Q(
        n624) );
  MUX21X1 U1668 ( .IN1(\regfile[13][14] ), .IN2(AluOut[14]), .S(n1289), .Q(
        n623) );
  MUX21X1 U1669 ( .IN1(\regfile[14][14] ), .IN2(AluOut[14]), .S(n1290), .Q(
        n622) );
  MUX21X1 U1670 ( .IN1(\regfile[15][14] ), .IN2(AluOut[14]), .S(n1291), .Q(
        n621) );
  AO221X1 U1671 ( .IN1(n1268), .IN2(AluOut[13]), .IN3(N236), .IN4(n1269), 
        .IN5(n1360), .Q(n620) );
  AO21X1 U1672 ( .IN1(n1008), .IN2(IFID_A[13]), .IN3(n1361), .Q(n1360) );
  MUX21X1 U1673 ( .IN1(n1362), .IN2(n1363), .S(IFID_B[13]), .Q(n1361) );
  AO21X1 U1674 ( .IN1(n1274), .IN2(IFID_A[13]), .IN3(n1009), .Q(n1363) );
  NOR2X0 U1675 ( .IN1(n1275), .IN2(IFID_A[13]), .QN(n1362) );
  MUX21X1 U1676 ( .IN1(\regfile[0][13] ), .IN2(AluOut[13]), .S(n1276), .Q(n619) );
  MUX21X1 U1677 ( .IN1(\regfile[1][13] ), .IN2(AluOut[13]), .S(n1277), .Q(n618) );
  MUX21X1 U1678 ( .IN1(\regfile[2][13] ), .IN2(AluOut[13]), .S(n1278), .Q(n617) );
  MUX21X1 U1679 ( .IN1(\regfile[3][13] ), .IN2(AluOut[13]), .S(n1279), .Q(n616) );
  MUX21X1 U1680 ( .IN1(\regfile[4][13] ), .IN2(AluOut[13]), .S(n1280), .Q(n615) );
  MUX21X1 U1681 ( .IN1(\regfile[5][13] ), .IN2(AluOut[13]), .S(n1281), .Q(n614) );
  MUX21X1 U1682 ( .IN1(\regfile[6][13] ), .IN2(AluOut[13]), .S(n1282), .Q(n613) );
  MUX21X1 U1683 ( .IN1(\regfile[7][13] ), .IN2(AluOut[13]), .S(n1283), .Q(n612) );
  MUX21X1 U1684 ( .IN1(\regfile[8][13] ), .IN2(AluOut[13]), .S(n1284), .Q(n611) );
  MUX21X1 U1685 ( .IN1(\regfile[9][13] ), .IN2(AluOut[13]), .S(n1285), .Q(n610) );
  MUX21X1 U1686 ( .IN1(\regfile[10][13] ), .IN2(AluOut[13]), .S(n1286), .Q(
        n609) );
  MUX21X1 U1687 ( .IN1(\regfile[11][13] ), .IN2(AluOut[13]), .S(n1287), .Q(
        n608) );
  MUX21X1 U1688 ( .IN1(\regfile[12][13] ), .IN2(AluOut[13]), .S(n1288), .Q(
        n607) );
  MUX21X1 U1689 ( .IN1(\regfile[13][13] ), .IN2(AluOut[13]), .S(n1289), .Q(
        n606) );
  MUX21X1 U1690 ( .IN1(\regfile[14][13] ), .IN2(AluOut[13]), .S(n1290), .Q(
        n605) );
  MUX21X1 U1691 ( .IN1(\regfile[15][13] ), .IN2(AluOut[13]), .S(n1291), .Q(
        n604) );
  AO221X1 U1692 ( .IN1(n1268), .IN2(AluOut[12]), .IN3(N235), .IN4(n1269), 
        .IN5(n1364), .Q(n603) );
  AO21X1 U1693 ( .IN1(n1011), .IN2(IFID_A[12]), .IN3(n1365), .Q(n1364) );
  MUX21X1 U1694 ( .IN1(n1366), .IN2(n1367), .S(IFID_B[12]), .Q(n1365) );
  AO21X1 U1695 ( .IN1(n1274), .IN2(IFID_A[12]), .IN3(n1008), .Q(n1367) );
  NOR2X0 U1696 ( .IN1(n1275), .IN2(IFID_A[12]), .QN(n1366) );
  MUX21X1 U1697 ( .IN1(\regfile[0][12] ), .IN2(AluOut[12]), .S(n1276), .Q(n602) );
  MUX21X1 U1698 ( .IN1(\regfile[1][12] ), .IN2(AluOut[12]), .S(n1277), .Q(n601) );
  MUX21X1 U1699 ( .IN1(\regfile[2][12] ), .IN2(AluOut[12]), .S(n1278), .Q(n600) );
  MUX21X1 U1700 ( .IN1(\regfile[3][12] ), .IN2(AluOut[12]), .S(n1279), .Q(n599) );
  MUX21X1 U1701 ( .IN1(\regfile[4][12] ), .IN2(AluOut[12]), .S(n1280), .Q(n598) );
  MUX21X1 U1702 ( .IN1(\regfile[5][12] ), .IN2(AluOut[12]), .S(n1281), .Q(n597) );
  MUX21X1 U1703 ( .IN1(\regfile[6][12] ), .IN2(AluOut[12]), .S(n1282), .Q(n596) );
  MUX21X1 U1704 ( .IN1(\regfile[7][12] ), .IN2(AluOut[12]), .S(n1283), .Q(n595) );
  MUX21X1 U1705 ( .IN1(\regfile[8][12] ), .IN2(AluOut[12]), .S(n1284), .Q(n594) );
  MUX21X1 U1706 ( .IN1(\regfile[9][12] ), .IN2(AluOut[12]), .S(n1285), .Q(n593) );
  MUX21X1 U1707 ( .IN1(\regfile[10][12] ), .IN2(AluOut[12]), .S(n1286), .Q(
        n592) );
  MUX21X1 U1708 ( .IN1(\regfile[11][12] ), .IN2(AluOut[12]), .S(n1287), .Q(
        n591) );
  MUX21X1 U1709 ( .IN1(\regfile[12][12] ), .IN2(AluOut[12]), .S(n1288), .Q(
        n590) );
  MUX21X1 U1710 ( .IN1(\regfile[13][12] ), .IN2(AluOut[12]), .S(n1289), .Q(
        n589) );
  MUX21X1 U1711 ( .IN1(\regfile[14][12] ), .IN2(AluOut[12]), .S(n1290), .Q(
        n588) );
  MUX21X1 U1712 ( .IN1(\regfile[15][12] ), .IN2(AluOut[12]), .S(n1291), .Q(
        n587) );
  AO221X1 U1713 ( .IN1(n1268), .IN2(AluOut[11]), .IN3(N234), .IN4(n1269), 
        .IN5(n1368), .Q(n586) );
  AO21X1 U1714 ( .IN1(n1010), .IN2(IFID_A[11]), .IN3(n1369), .Q(n1368) );
  MUX21X1 U1715 ( .IN1(n1370), .IN2(n1371), .S(IFID_B[11]), .Q(n1369) );
  AO21X1 U1716 ( .IN1(n1274), .IN2(IFID_A[11]), .IN3(n1011), .Q(n1371) );
  NOR2X0 U1717 ( .IN1(n1275), .IN2(IFID_A[11]), .QN(n1370) );
  MUX21X1 U1718 ( .IN1(\regfile[0][11] ), .IN2(AluOut[11]), .S(n1276), .Q(n585) );
  MUX21X1 U1719 ( .IN1(\regfile[1][11] ), .IN2(AluOut[11]), .S(n1277), .Q(n584) );
  MUX21X1 U1720 ( .IN1(\regfile[2][11] ), .IN2(AluOut[11]), .S(n1278), .Q(n583) );
  MUX21X1 U1721 ( .IN1(\regfile[3][11] ), .IN2(AluOut[11]), .S(n1279), .Q(n582) );
  MUX21X1 U1722 ( .IN1(\regfile[4][11] ), .IN2(AluOut[11]), .S(n1280), .Q(n581) );
  MUX21X1 U1723 ( .IN1(\regfile[5][11] ), .IN2(AluOut[11]), .S(n1281), .Q(n580) );
  MUX21X1 U1724 ( .IN1(\regfile[6][11] ), .IN2(AluOut[11]), .S(n1282), .Q(n579) );
  MUX21X1 U1725 ( .IN1(\regfile[7][11] ), .IN2(AluOut[11]), .S(n1283), .Q(n578) );
  MUX21X1 U1726 ( .IN1(\regfile[8][11] ), .IN2(AluOut[11]), .S(n1284), .Q(n577) );
  MUX21X1 U1727 ( .IN1(\regfile[9][11] ), .IN2(AluOut[11]), .S(n1285), .Q(n576) );
  MUX21X1 U1728 ( .IN1(\regfile[10][11] ), .IN2(AluOut[11]), .S(n1286), .Q(
        n575) );
  MUX21X1 U1729 ( .IN1(\regfile[11][11] ), .IN2(AluOut[11]), .S(n1287), .Q(
        n574) );
  MUX21X1 U1730 ( .IN1(\regfile[12][11] ), .IN2(AluOut[11]), .S(n1288), .Q(
        n573) );
  MUX21X1 U1731 ( .IN1(\regfile[13][11] ), .IN2(AluOut[11]), .S(n1289), .Q(
        n572) );
  MUX21X1 U1732 ( .IN1(\regfile[14][11] ), .IN2(AluOut[11]), .S(n1290), .Q(
        n571) );
  MUX21X1 U1733 ( .IN1(\regfile[15][11] ), .IN2(AluOut[11]), .S(n1291), .Q(
        n570) );
  AO221X1 U1734 ( .IN1(n1268), .IN2(AluOut[10]), .IN3(N233), .IN4(n1269), 
        .IN5(n1372), .Q(n569) );
  AO21X1 U1735 ( .IN1(n1009), .IN2(IFID_A[10]), .IN3(n1373), .Q(n1372) );
  MUX21X1 U1736 ( .IN1(n1374), .IN2(n1375), .S(IFID_B[10]), .Q(n1373) );
  AO21X1 U1737 ( .IN1(n1274), .IN2(IFID_A[10]), .IN3(n1010), .Q(n1375) );
  NOR2X0 U1738 ( .IN1(n1275), .IN2(IFID_A[10]), .QN(n1374) );
  MUX21X1 U1739 ( .IN1(\regfile[0][10] ), .IN2(AluOut[10]), .S(n1276), .Q(n568) );
  MUX21X1 U1740 ( .IN1(\regfile[1][10] ), .IN2(AluOut[10]), .S(n1277), .Q(n567) );
  MUX21X1 U1741 ( .IN1(\regfile[2][10] ), .IN2(AluOut[10]), .S(n1278), .Q(n566) );
  MUX21X1 U1742 ( .IN1(\regfile[3][10] ), .IN2(AluOut[10]), .S(n1279), .Q(n565) );
  MUX21X1 U1743 ( .IN1(\regfile[4][10] ), .IN2(AluOut[10]), .S(n1280), .Q(n564) );
  MUX21X1 U1744 ( .IN1(\regfile[5][10] ), .IN2(AluOut[10]), .S(n1281), .Q(n563) );
  MUX21X1 U1745 ( .IN1(\regfile[6][10] ), .IN2(AluOut[10]), .S(n1282), .Q(n562) );
  MUX21X1 U1746 ( .IN1(\regfile[7][10] ), .IN2(AluOut[10]), .S(n1283), .Q(n561) );
  MUX21X1 U1747 ( .IN1(\regfile[8][10] ), .IN2(AluOut[10]), .S(n1284), .Q(n560) );
  MUX21X1 U1748 ( .IN1(\regfile[9][10] ), .IN2(AluOut[10]), .S(n1285), .Q(n559) );
  MUX21X1 U1749 ( .IN1(\regfile[10][10] ), .IN2(AluOut[10]), .S(n1286), .Q(
        n558) );
  MUX21X1 U1750 ( .IN1(\regfile[11][10] ), .IN2(AluOut[10]), .S(n1287), .Q(
        n557) );
  MUX21X1 U1751 ( .IN1(\regfile[12][10] ), .IN2(AluOut[10]), .S(n1288), .Q(
        n556) );
  MUX21X1 U1752 ( .IN1(\regfile[13][10] ), .IN2(AluOut[10]), .S(n1289), .Q(
        n555) );
  MUX21X1 U1753 ( .IN1(\regfile[14][10] ), .IN2(AluOut[10]), .S(n1290), .Q(
        n554) );
  MUX21X1 U1754 ( .IN1(\regfile[15][10] ), .IN2(AluOut[10]), .S(n1291), .Q(
        n553) );
  AO221X1 U1755 ( .IN1(n1268), .IN2(AluOut[9]), .IN3(N232), .IN4(n1269), .IN5(
        n1376), .Q(n552) );
  AO21X1 U1756 ( .IN1(n1008), .IN2(IFID_A[9]), .IN3(n1377), .Q(n1376) );
  MUX21X1 U1757 ( .IN1(n1378), .IN2(n1379), .S(IFID_B[9]), .Q(n1377) );
  AO21X1 U1758 ( .IN1(n1274), .IN2(IFID_A[9]), .IN3(n1009), .Q(n1379) );
  NOR2X0 U1759 ( .IN1(n1275), .IN2(IFID_A[9]), .QN(n1378) );
  MUX21X1 U1760 ( .IN1(\regfile[0][9] ), .IN2(AluOut[9]), .S(n1276), .Q(n551)
         );
  MUX21X1 U1761 ( .IN1(\regfile[1][9] ), .IN2(AluOut[9]), .S(n1277), .Q(n550)
         );
  MUX21X1 U1762 ( .IN1(\regfile[2][9] ), .IN2(AluOut[9]), .S(n1278), .Q(n549)
         );
  MUX21X1 U1763 ( .IN1(\regfile[3][9] ), .IN2(AluOut[9]), .S(n1279), .Q(n548)
         );
  MUX21X1 U1764 ( .IN1(\regfile[4][9] ), .IN2(AluOut[9]), .S(n1280), .Q(n547)
         );
  MUX21X1 U1765 ( .IN1(\regfile[5][9] ), .IN2(AluOut[9]), .S(n1281), .Q(n546)
         );
  MUX21X1 U1766 ( .IN1(\regfile[6][9] ), .IN2(AluOut[9]), .S(n1282), .Q(n545)
         );
  MUX21X1 U1767 ( .IN1(\regfile[7][9] ), .IN2(AluOut[9]), .S(n1283), .Q(n544)
         );
  MUX21X1 U1768 ( .IN1(\regfile[8][9] ), .IN2(AluOut[9]), .S(n1284), .Q(n543)
         );
  MUX21X1 U1769 ( .IN1(\regfile[9][9] ), .IN2(AluOut[9]), .S(n1285), .Q(n542)
         );
  MUX21X1 U1770 ( .IN1(\regfile[10][9] ), .IN2(AluOut[9]), .S(n1286), .Q(n541)
         );
  MUX21X1 U1771 ( .IN1(\regfile[11][9] ), .IN2(AluOut[9]), .S(n1287), .Q(n540)
         );
  MUX21X1 U1772 ( .IN1(\regfile[12][9] ), .IN2(AluOut[9]), .S(n1288), .Q(n539)
         );
  MUX21X1 U1773 ( .IN1(\regfile[13][9] ), .IN2(AluOut[9]), .S(n1289), .Q(n538)
         );
  MUX21X1 U1774 ( .IN1(\regfile[14][9] ), .IN2(AluOut[9]), .S(n1290), .Q(n537)
         );
  MUX21X1 U1775 ( .IN1(\regfile[15][9] ), .IN2(AluOut[9]), .S(n1291), .Q(n536)
         );
  AO221X1 U1776 ( .IN1(n1268), .IN2(AluOut[8]), .IN3(N231), .IN4(n1269), .IN5(
        n1380), .Q(n535) );
  AO21X1 U1777 ( .IN1(n1011), .IN2(IFID_A[8]), .IN3(n1381), .Q(n1380) );
  MUX21X1 U1778 ( .IN1(n1382), .IN2(n1383), .S(IFID_B[8]), .Q(n1381) );
  AO21X1 U1779 ( .IN1(n1274), .IN2(IFID_A[8]), .IN3(n1008), .Q(n1383) );
  NOR2X0 U1780 ( .IN1(n1275), .IN2(IFID_A[8]), .QN(n1382) );
  MUX21X1 U1781 ( .IN1(\regfile[0][8] ), .IN2(AluOut[8]), .S(n1276), .Q(n534)
         );
  MUX21X1 U1782 ( .IN1(\regfile[1][8] ), .IN2(AluOut[8]), .S(n1277), .Q(n533)
         );
  MUX21X1 U1783 ( .IN1(\regfile[2][8] ), .IN2(AluOut[8]), .S(n1278), .Q(n532)
         );
  MUX21X1 U1784 ( .IN1(\regfile[3][8] ), .IN2(AluOut[8]), .S(n1279), .Q(n531)
         );
  MUX21X1 U1785 ( .IN1(\regfile[4][8] ), .IN2(AluOut[8]), .S(n1280), .Q(n530)
         );
  MUX21X1 U1786 ( .IN1(\regfile[5][8] ), .IN2(AluOut[8]), .S(n1281), .Q(n529)
         );
  MUX21X1 U1787 ( .IN1(\regfile[6][8] ), .IN2(AluOut[8]), .S(n1282), .Q(n528)
         );
  MUX21X1 U1788 ( .IN1(\regfile[7][8] ), .IN2(AluOut[8]), .S(n1283), .Q(n527)
         );
  MUX21X1 U1789 ( .IN1(\regfile[8][8] ), .IN2(AluOut[8]), .S(n1284), .Q(n526)
         );
  MUX21X1 U1790 ( .IN1(\regfile[9][8] ), .IN2(AluOut[8]), .S(n1285), .Q(n525)
         );
  MUX21X1 U1791 ( .IN1(\regfile[10][8] ), .IN2(AluOut[8]), .S(n1286), .Q(n524)
         );
  MUX21X1 U1792 ( .IN1(\regfile[11][8] ), .IN2(AluOut[8]), .S(n1287), .Q(n523)
         );
  MUX21X1 U1793 ( .IN1(\regfile[12][8] ), .IN2(AluOut[8]), .S(n1288), .Q(n522)
         );
  MUX21X1 U1794 ( .IN1(\regfile[13][8] ), .IN2(AluOut[8]), .S(n1289), .Q(n521)
         );
  MUX21X1 U1795 ( .IN1(\regfile[14][8] ), .IN2(AluOut[8]), .S(n1290), .Q(n520)
         );
  MUX21X1 U1796 ( .IN1(\regfile[15][8] ), .IN2(AluOut[8]), .S(n1291), .Q(n519)
         );
  AO221X1 U1797 ( .IN1(n1268), .IN2(AluOut[7]), .IN3(N230), .IN4(n1269), .IN5(
        n1384), .Q(n518) );
  AO21X1 U1798 ( .IN1(n1010), .IN2(IFID_A[7]), .IN3(n1385), .Q(n1384) );
  MUX21X1 U1799 ( .IN1(n1386), .IN2(n1387), .S(IFID_B[7]), .Q(n1385) );
  AO21X1 U1800 ( .IN1(n1274), .IN2(IFID_A[7]), .IN3(n1011), .Q(n1387) );
  NOR2X0 U1801 ( .IN1(n1275), .IN2(IFID_A[7]), .QN(n1386) );
  MUX21X1 U1802 ( .IN1(\regfile[0][7] ), .IN2(AluOut[7]), .S(n1276), .Q(n517)
         );
  MUX21X1 U1803 ( .IN1(\regfile[1][7] ), .IN2(AluOut[7]), .S(n1277), .Q(n516)
         );
  MUX21X1 U1804 ( .IN1(\regfile[2][7] ), .IN2(AluOut[7]), .S(n1278), .Q(n515)
         );
  MUX21X1 U1805 ( .IN1(\regfile[3][7] ), .IN2(AluOut[7]), .S(n1279), .Q(n514)
         );
  MUX21X1 U1806 ( .IN1(\regfile[4][7] ), .IN2(AluOut[7]), .S(n1280), .Q(n513)
         );
  MUX21X1 U1807 ( .IN1(\regfile[5][7] ), .IN2(AluOut[7]), .S(n1281), .Q(n512)
         );
  MUX21X1 U1808 ( .IN1(\regfile[6][7] ), .IN2(AluOut[7]), .S(n1282), .Q(n511)
         );
  MUX21X1 U1809 ( .IN1(\regfile[7][7] ), .IN2(AluOut[7]), .S(n1283), .Q(n510)
         );
  MUX21X1 U1810 ( .IN1(\regfile[8][7] ), .IN2(AluOut[7]), .S(n1284), .Q(n509)
         );
  MUX21X1 U1811 ( .IN1(\regfile[9][7] ), .IN2(AluOut[7]), .S(n1285), .Q(n508)
         );
  MUX21X1 U1812 ( .IN1(\regfile[10][7] ), .IN2(AluOut[7]), .S(n1286), .Q(n507)
         );
  MUX21X1 U1813 ( .IN1(\regfile[11][7] ), .IN2(AluOut[7]), .S(n1287), .Q(n506)
         );
  MUX21X1 U1814 ( .IN1(\regfile[12][7] ), .IN2(AluOut[7]), .S(n1288), .Q(n505)
         );
  MUX21X1 U1815 ( .IN1(\regfile[13][7] ), .IN2(AluOut[7]), .S(n1289), .Q(n504)
         );
  MUX21X1 U1816 ( .IN1(\regfile[14][7] ), .IN2(AluOut[7]), .S(n1290), .Q(n503)
         );
  MUX21X1 U1817 ( .IN1(\regfile[15][7] ), .IN2(AluOut[7]), .S(n1291), .Q(n502)
         );
  AO221X1 U1818 ( .IN1(n1268), .IN2(AluOut[6]), .IN3(N229), .IN4(n1269), .IN5(
        n1388), .Q(n501) );
  AO21X1 U1819 ( .IN1(n1009), .IN2(IFID_A[6]), .IN3(n1389), .Q(n1388) );
  MUX21X1 U1820 ( .IN1(n1390), .IN2(n1391), .S(IFID_B[6]), .Q(n1389) );
  AO21X1 U1821 ( .IN1(n1274), .IN2(IFID_A[6]), .IN3(n1010), .Q(n1391) );
  NOR2X0 U1822 ( .IN1(n1275), .IN2(IFID_A[6]), .QN(n1390) );
  MUX21X1 U1823 ( .IN1(\regfile[0][6] ), .IN2(AluOut[6]), .S(n1276), .Q(n500)
         );
  MUX21X1 U1824 ( .IN1(\regfile[1][6] ), .IN2(AluOut[6]), .S(n1277), .Q(n499)
         );
  MUX21X1 U1825 ( .IN1(\regfile[2][6] ), .IN2(AluOut[6]), .S(n1278), .Q(n498)
         );
  MUX21X1 U1826 ( .IN1(\regfile[3][6] ), .IN2(AluOut[6]), .S(n1279), .Q(n497)
         );
  MUX21X1 U1827 ( .IN1(\regfile[4][6] ), .IN2(AluOut[6]), .S(n1280), .Q(n496)
         );
  MUX21X1 U1828 ( .IN1(\regfile[5][6] ), .IN2(AluOut[6]), .S(n1281), .Q(n495)
         );
  MUX21X1 U1829 ( .IN1(\regfile[6][6] ), .IN2(AluOut[6]), .S(n1282), .Q(n494)
         );
  MUX21X1 U1830 ( .IN1(\regfile[7][6] ), .IN2(AluOut[6]), .S(n1283), .Q(n493)
         );
  MUX21X1 U1831 ( .IN1(\regfile[8][6] ), .IN2(AluOut[6]), .S(n1284), .Q(n492)
         );
  MUX21X1 U1832 ( .IN1(\regfile[9][6] ), .IN2(AluOut[6]), .S(n1285), .Q(n491)
         );
  MUX21X1 U1833 ( .IN1(\regfile[10][6] ), .IN2(AluOut[6]), .S(n1286), .Q(n490)
         );
  MUX21X1 U1834 ( .IN1(\regfile[11][6] ), .IN2(AluOut[6]), .S(n1287), .Q(n489)
         );
  MUX21X1 U1835 ( .IN1(\regfile[12][6] ), .IN2(AluOut[6]), .S(n1288), .Q(n488)
         );
  MUX21X1 U1836 ( .IN1(\regfile[13][6] ), .IN2(AluOut[6]), .S(n1289), .Q(n487)
         );
  MUX21X1 U1837 ( .IN1(\regfile[14][6] ), .IN2(AluOut[6]), .S(n1290), .Q(n486)
         );
  MUX21X1 U1838 ( .IN1(\regfile[15][6] ), .IN2(AluOut[6]), .S(n1291), .Q(n485)
         );
  AO221X1 U1839 ( .IN1(n1268), .IN2(AluOut[5]), .IN3(N228), .IN4(n1269), .IN5(
        n1392), .Q(n484) );
  AO21X1 U1840 ( .IN1(n1008), .IN2(IFID_A[5]), .IN3(n1393), .Q(n1392) );
  MUX21X1 U1841 ( .IN1(n1394), .IN2(n1395), .S(IFID_B[5]), .Q(n1393) );
  AO21X1 U1842 ( .IN1(n1274), .IN2(IFID_A[5]), .IN3(n1009), .Q(n1395) );
  NOR2X0 U1843 ( .IN1(n1275), .IN2(IFID_A[5]), .QN(n1394) );
  MUX21X1 U1844 ( .IN1(\regfile[0][5] ), .IN2(AluOut[5]), .S(n1276), .Q(n483)
         );
  MUX21X1 U1845 ( .IN1(\regfile[1][5] ), .IN2(AluOut[5]), .S(n1277), .Q(n482)
         );
  MUX21X1 U1846 ( .IN1(\regfile[2][5] ), .IN2(AluOut[5]), .S(n1278), .Q(n481)
         );
  MUX21X1 U1847 ( .IN1(\regfile[3][5] ), .IN2(AluOut[5]), .S(n1279), .Q(n480)
         );
  MUX21X1 U1848 ( .IN1(\regfile[4][5] ), .IN2(AluOut[5]), .S(n1280), .Q(n479)
         );
  MUX21X1 U1849 ( .IN1(\regfile[5][5] ), .IN2(AluOut[5]), .S(n1281), .Q(n478)
         );
  MUX21X1 U1850 ( .IN1(\regfile[6][5] ), .IN2(AluOut[5]), .S(n1282), .Q(n477)
         );
  MUX21X1 U1851 ( .IN1(\regfile[7][5] ), .IN2(AluOut[5]), .S(n1283), .Q(n476)
         );
  MUX21X1 U1852 ( .IN1(\regfile[8][5] ), .IN2(AluOut[5]), .S(n1284), .Q(n475)
         );
  MUX21X1 U1853 ( .IN1(\regfile[9][5] ), .IN2(AluOut[5]), .S(n1285), .Q(n474)
         );
  MUX21X1 U1854 ( .IN1(\regfile[10][5] ), .IN2(AluOut[5]), .S(n1286), .Q(n473)
         );
  MUX21X1 U1855 ( .IN1(\regfile[11][5] ), .IN2(AluOut[5]), .S(n1287), .Q(n472)
         );
  MUX21X1 U1856 ( .IN1(\regfile[12][5] ), .IN2(AluOut[5]), .S(n1288), .Q(n471)
         );
  MUX21X1 U1857 ( .IN1(\regfile[13][5] ), .IN2(AluOut[5]), .S(n1289), .Q(n470)
         );
  MUX21X1 U1858 ( .IN1(\regfile[14][5] ), .IN2(AluOut[5]), .S(n1290), .Q(n469)
         );
  MUX21X1 U1859 ( .IN1(\regfile[15][5] ), .IN2(AluOut[5]), .S(n1291), .Q(n468)
         );
  AO221X1 U1860 ( .IN1(n1268), .IN2(AluOut[4]), .IN3(N227), .IN4(n1269), .IN5(
        n1396), .Q(n467) );
  AO21X1 U1861 ( .IN1(n1011), .IN2(IFID_A[4]), .IN3(n1397), .Q(n1396) );
  MUX21X1 U1862 ( .IN1(n1398), .IN2(n1399), .S(IFID_B[4]), .Q(n1397) );
  AO21X1 U1863 ( .IN1(n1274), .IN2(IFID_A[4]), .IN3(n1008), .Q(n1399) );
  NOR2X0 U1864 ( .IN1(n1275), .IN2(IFID_A[4]), .QN(n1398) );
  MUX21X1 U1865 ( .IN1(\regfile[0][4] ), .IN2(AluOut[4]), .S(n1276), .Q(n466)
         );
  MUX21X1 U1866 ( .IN1(\regfile[1][4] ), .IN2(AluOut[4]), .S(n1277), .Q(n465)
         );
  MUX21X1 U1867 ( .IN1(\regfile[2][4] ), .IN2(AluOut[4]), .S(n1278), .Q(n464)
         );
  MUX21X1 U1868 ( .IN1(\regfile[3][4] ), .IN2(AluOut[4]), .S(n1279), .Q(n463)
         );
  MUX21X1 U1869 ( .IN1(\regfile[4][4] ), .IN2(AluOut[4]), .S(n1280), .Q(n462)
         );
  MUX21X1 U1870 ( .IN1(\regfile[5][4] ), .IN2(AluOut[4]), .S(n1281), .Q(n461)
         );
  MUX21X1 U1871 ( .IN1(\regfile[6][4] ), .IN2(AluOut[4]), .S(n1282), .Q(n460)
         );
  MUX21X1 U1872 ( .IN1(\regfile[7][4] ), .IN2(AluOut[4]), .S(n1283), .Q(n459)
         );
  MUX21X1 U1873 ( .IN1(\regfile[8][4] ), .IN2(AluOut[4]), .S(n1284), .Q(n458)
         );
  MUX21X1 U1874 ( .IN1(\regfile[9][4] ), .IN2(AluOut[4]), .S(n1285), .Q(n457)
         );
  MUX21X1 U1875 ( .IN1(\regfile[10][4] ), .IN2(AluOut[4]), .S(n1286), .Q(n456)
         );
  MUX21X1 U1876 ( .IN1(\regfile[11][4] ), .IN2(AluOut[4]), .S(n1287), .Q(n455)
         );
  MUX21X1 U1877 ( .IN1(\regfile[12][4] ), .IN2(AluOut[4]), .S(n1288), .Q(n454)
         );
  MUX21X1 U1878 ( .IN1(\regfile[13][4] ), .IN2(AluOut[4]), .S(n1289), .Q(n453)
         );
  MUX21X1 U1879 ( .IN1(\regfile[14][4] ), .IN2(AluOut[4]), .S(n1290), .Q(n452)
         );
  MUX21X1 U1880 ( .IN1(\regfile[15][4] ), .IN2(AluOut[4]), .S(n1291), .Q(n451)
         );
  AO221X1 U1881 ( .IN1(n1268), .IN2(AluOut[3]), .IN3(N226), .IN4(n1269), .IN5(
        n1400), .Q(n450) );
  AO21X1 U1882 ( .IN1(n1010), .IN2(IFID_A[3]), .IN3(n1401), .Q(n1400) );
  MUX21X1 U1883 ( .IN1(n1402), .IN2(n1403), .S(IFID_B[3]), .Q(n1401) );
  AO21X1 U1884 ( .IN1(n1274), .IN2(IFID_A[3]), .IN3(n1011), .Q(n1403) );
  NOR2X0 U1885 ( .IN1(n1275), .IN2(IFID_A[3]), .QN(n1402) );
  MUX21X1 U1886 ( .IN1(\regfile[0][3] ), .IN2(AluOut[3]), .S(n1276), .Q(n449)
         );
  MUX21X1 U1887 ( .IN1(\regfile[1][3] ), .IN2(AluOut[3]), .S(n1277), .Q(n448)
         );
  MUX21X1 U1888 ( .IN1(\regfile[2][3] ), .IN2(AluOut[3]), .S(n1278), .Q(n447)
         );
  MUX21X1 U1889 ( .IN1(\regfile[3][3] ), .IN2(AluOut[3]), .S(n1279), .Q(n446)
         );
  MUX21X1 U1890 ( .IN1(\regfile[4][3] ), .IN2(AluOut[3]), .S(n1280), .Q(n445)
         );
  MUX21X1 U1891 ( .IN1(\regfile[5][3] ), .IN2(AluOut[3]), .S(n1281), .Q(n444)
         );
  MUX21X1 U1892 ( .IN1(\regfile[6][3] ), .IN2(AluOut[3]), .S(n1282), .Q(n443)
         );
  MUX21X1 U1893 ( .IN1(\regfile[7][3] ), .IN2(AluOut[3]), .S(n1283), .Q(n442)
         );
  MUX21X1 U1894 ( .IN1(\regfile[8][3] ), .IN2(AluOut[3]), .S(n1284), .Q(n441)
         );
  MUX21X1 U1895 ( .IN1(\regfile[9][3] ), .IN2(AluOut[3]), .S(n1285), .Q(n440)
         );
  MUX21X1 U1896 ( .IN1(\regfile[10][3] ), .IN2(AluOut[3]), .S(n1286), .Q(n439)
         );
  MUX21X1 U1897 ( .IN1(\regfile[11][3] ), .IN2(AluOut[3]), .S(n1287), .Q(n438)
         );
  MUX21X1 U1898 ( .IN1(\regfile[12][3] ), .IN2(AluOut[3]), .S(n1288), .Q(n437)
         );
  MUX21X1 U1899 ( .IN1(\regfile[13][3] ), .IN2(AluOut[3]), .S(n1289), .Q(n436)
         );
  MUX21X1 U1900 ( .IN1(\regfile[14][3] ), .IN2(AluOut[3]), .S(n1290), .Q(n435)
         );
  MUX21X1 U1901 ( .IN1(\regfile[15][3] ), .IN2(AluOut[3]), .S(n1291), .Q(n434)
         );
  AO221X1 U1902 ( .IN1(n1268), .IN2(AluOut[2]), .IN3(N225), .IN4(n1269), .IN5(
        n1404), .Q(n433) );
  AO21X1 U1903 ( .IN1(n1009), .IN2(IFID_A[2]), .IN3(n1405), .Q(n1404) );
  MUX21X1 U1904 ( .IN1(n1406), .IN2(n1407), .S(IFID_B[2]), .Q(n1405) );
  AO21X1 U1905 ( .IN1(n1274), .IN2(IFID_A[2]), .IN3(n1010), .Q(n1407) );
  NOR2X0 U1906 ( .IN1(n1275), .IN2(IFID_A[2]), .QN(n1406) );
  MUX21X1 U1907 ( .IN1(\regfile[0][2] ), .IN2(AluOut[2]), .S(n1276), .Q(n432)
         );
  MUX21X1 U1908 ( .IN1(\regfile[1][2] ), .IN2(AluOut[2]), .S(n1277), .Q(n431)
         );
  MUX21X1 U1909 ( .IN1(\regfile[2][2] ), .IN2(AluOut[2]), .S(n1278), .Q(n430)
         );
  MUX21X1 U1910 ( .IN1(\regfile[3][2] ), .IN2(AluOut[2]), .S(n1279), .Q(n429)
         );
  MUX21X1 U1911 ( .IN1(\regfile[4][2] ), .IN2(AluOut[2]), .S(n1280), .Q(n428)
         );
  MUX21X1 U1912 ( .IN1(\regfile[5][2] ), .IN2(AluOut[2]), .S(n1281), .Q(n427)
         );
  MUX21X1 U1913 ( .IN1(\regfile[6][2] ), .IN2(AluOut[2]), .S(n1282), .Q(n426)
         );
  MUX21X1 U1914 ( .IN1(\regfile[7][2] ), .IN2(AluOut[2]), .S(n1283), .Q(n425)
         );
  MUX21X1 U1915 ( .IN1(\regfile[8][2] ), .IN2(AluOut[2]), .S(n1284), .Q(n424)
         );
  MUX21X1 U1916 ( .IN1(\regfile[9][2] ), .IN2(AluOut[2]), .S(n1285), .Q(n423)
         );
  MUX21X1 U1917 ( .IN1(\regfile[10][2] ), .IN2(AluOut[2]), .S(n1286), .Q(n422)
         );
  MUX21X1 U1918 ( .IN1(\regfile[11][2] ), .IN2(AluOut[2]), .S(n1287), .Q(n421)
         );
  MUX21X1 U1919 ( .IN1(\regfile[12][2] ), .IN2(AluOut[2]), .S(n1288), .Q(n420)
         );
  MUX21X1 U1920 ( .IN1(\regfile[13][2] ), .IN2(AluOut[2]), .S(n1289), .Q(n419)
         );
  MUX21X1 U1921 ( .IN1(\regfile[14][2] ), .IN2(AluOut[2]), .S(n1290), .Q(n418)
         );
  MUX21X1 U1922 ( .IN1(\regfile[15][2] ), .IN2(AluOut[2]), .S(n1291), .Q(n417)
         );
  AO221X1 U1923 ( .IN1(n1268), .IN2(AluOut[1]), .IN3(N224), .IN4(n1269), .IN5(
        n1408), .Q(n416) );
  AO21X1 U1924 ( .IN1(n1008), .IN2(IFID_A[1]), .IN3(n1409), .Q(n1408) );
  MUX21X1 U1925 ( .IN1(n1410), .IN2(n1411), .S(IFID_B[1]), .Q(n1409) );
  AO21X1 U1926 ( .IN1(n1274), .IN2(IFID_A[1]), .IN3(n1009), .Q(n1411) );
  NOR2X0 U1927 ( .IN1(n1275), .IN2(IFID_A[1]), .QN(n1410) );
  INVX0 U1928 ( .INP(n1412), .ZN(n1268) );
  MUX21X1 U1929 ( .IN1(\regfile[0][1] ), .IN2(AluOut[1]), .S(n1276), .Q(n415)
         );
  MUX21X1 U1930 ( .IN1(\regfile[1][1] ), .IN2(AluOut[1]), .S(n1277), .Q(n414)
         );
  MUX21X1 U1931 ( .IN1(\regfile[2][1] ), .IN2(AluOut[1]), .S(n1278), .Q(n413)
         );
  MUX21X1 U1932 ( .IN1(\regfile[3][1] ), .IN2(AluOut[1]), .S(n1279), .Q(n412)
         );
  MUX21X1 U1933 ( .IN1(\regfile[4][1] ), .IN2(AluOut[1]), .S(n1280), .Q(n411)
         );
  MUX21X1 U1934 ( .IN1(\regfile[5][1] ), .IN2(AluOut[1]), .S(n1281), .Q(n410)
         );
  MUX21X1 U1935 ( .IN1(\regfile[6][1] ), .IN2(AluOut[1]), .S(n1282), .Q(n409)
         );
  MUX21X1 U1936 ( .IN1(\regfile[7][1] ), .IN2(AluOut[1]), .S(n1283), .Q(n408)
         );
  MUX21X1 U1937 ( .IN1(\regfile[8][1] ), .IN2(AluOut[1]), .S(n1284), .Q(n407)
         );
  MUX21X1 U1938 ( .IN1(\regfile[9][1] ), .IN2(AluOut[1]), .S(n1285), .Q(n406)
         );
  MUX21X1 U1939 ( .IN1(\regfile[10][1] ), .IN2(AluOut[1]), .S(n1286), .Q(n405)
         );
  MUX21X1 U1940 ( .IN1(\regfile[11][1] ), .IN2(AluOut[1]), .S(n1287), .Q(n404)
         );
  MUX21X1 U1941 ( .IN1(\regfile[12][1] ), .IN2(AluOut[1]), .S(n1288), .Q(n403)
         );
  MUX21X1 U1942 ( .IN1(\regfile[13][1] ), .IN2(AluOut[1]), .S(n1289), .Q(n402)
         );
  MUX21X1 U1943 ( .IN1(\regfile[14][1] ), .IN2(AluOut[1]), .S(n1290), .Q(n401)
         );
  MUX21X1 U1944 ( .IN1(\regfile[15][1] ), .IN2(AluOut[1]), .S(n1291), .Q(n400)
         );
  NAND4X0 U1945 ( .IN1(n1413), .IN2(n1414), .IN3(n1415), .IN4(n1416), .QN(n399) );
  OA221X1 U1946 ( .IN1(n279), .IN2(n1412), .IN3(IFID_A[31]), .IN4(n1417), 
        .IN5(n1418), .Q(n1416) );
  AO22X1 U1947 ( .IN1(n1419), .IN2(n1420), .IN3(n1417), .IN4(n1421), .Q(n1418)
         );
  NAND3X0 U1948 ( .IN1(n346), .IN2(n1485), .IN3(n1422), .QN(n1421) );
  AO221X1 U1949 ( .IN1(n381), .IN2(IFID_A[30]), .IN3(n380), .IN4(IFID_A[29]), 
        .IN5(n1423), .Q(n1420) );
  OA221X1 U1950 ( .IN1(n380), .IN2(IFID_A[29]), .IN3(n379), .IN4(IFID_A[28]), 
        .IN5(n1424), .Q(n1423) );
  AO221X1 U1951 ( .IN1(n379), .IN2(IFID_A[28]), .IN3(n378), .IN4(IFID_A[27]), 
        .IN5(n1425), .Q(n1424) );
  OA221X1 U1952 ( .IN1(n378), .IN2(IFID_A[27]), .IN3(n377), .IN4(IFID_A[26]), 
        .IN5(n1426), .Q(n1425) );
  AO221X1 U1953 ( .IN1(n377), .IN2(IFID_A[26]), .IN3(n376), .IN4(IFID_A[25]), 
        .IN5(n1427), .Q(n1426) );
  OA221X1 U1954 ( .IN1(n376), .IN2(IFID_A[25]), .IN3(n375), .IN4(IFID_A[24]), 
        .IN5(n1428), .Q(n1427) );
  AO221X1 U1955 ( .IN1(n375), .IN2(IFID_A[24]), .IN3(n374), .IN4(IFID_A[23]), 
        .IN5(n1429), .Q(n1428) );
  OA221X1 U1956 ( .IN1(n374), .IN2(IFID_A[23]), .IN3(n373), .IN4(IFID_A[22]), 
        .IN5(n1430), .Q(n1429) );
  AO221X1 U1957 ( .IN1(n373), .IN2(IFID_A[22]), .IN3(n372), .IN4(IFID_A[21]), 
        .IN5(n1431), .Q(n1430) );
  OA221X1 U1958 ( .IN1(n372), .IN2(IFID_A[21]), .IN3(n371), .IN4(IFID_A[20]), 
        .IN5(n1432), .Q(n1431) );
  AO221X1 U1959 ( .IN1(n371), .IN2(IFID_A[20]), .IN3(n370), .IN4(IFID_A[19]), 
        .IN5(n1433), .Q(n1432) );
  OA221X1 U1960 ( .IN1(n370), .IN2(IFID_A[19]), .IN3(n369), .IN4(IFID_A[18]), 
        .IN5(n1434), .Q(n1433) );
  AO221X1 U1961 ( .IN1(n369), .IN2(IFID_A[18]), .IN3(n368), .IN4(IFID_A[17]), 
        .IN5(n1435), .Q(n1434) );
  OA221X1 U1962 ( .IN1(n368), .IN2(IFID_A[17]), .IN3(n367), .IN4(IFID_A[16]), 
        .IN5(n1436), .Q(n1435) );
  AO221X1 U1963 ( .IN1(n367), .IN2(IFID_A[16]), .IN3(n366), .IN4(IFID_A[15]), 
        .IN5(n1437), .Q(n1436) );
  OA221X1 U1964 ( .IN1(n366), .IN2(IFID_A[15]), .IN3(n365), .IN4(IFID_A[14]), 
        .IN5(n1438), .Q(n1437) );
  AO221X1 U1965 ( .IN1(n365), .IN2(IFID_A[14]), .IN3(n364), .IN4(IFID_A[13]), 
        .IN5(n1439), .Q(n1438) );
  OA221X1 U1966 ( .IN1(n364), .IN2(IFID_A[13]), .IN3(n363), .IN4(IFID_A[12]), 
        .IN5(n1440), .Q(n1439) );
  AO221X1 U1967 ( .IN1(n363), .IN2(IFID_A[12]), .IN3(n362), .IN4(IFID_A[11]), 
        .IN5(n1441), .Q(n1440) );
  OA221X1 U1968 ( .IN1(n362), .IN2(IFID_A[11]), .IN3(n361), .IN4(IFID_A[10]), 
        .IN5(n1442), .Q(n1441) );
  AO221X1 U1969 ( .IN1(n361), .IN2(IFID_A[10]), .IN3(n360), .IN4(IFID_A[9]), 
        .IN5(n1443), .Q(n1442) );
  OA221X1 U1970 ( .IN1(n360), .IN2(IFID_A[9]), .IN3(n359), .IN4(IFID_A[8]), 
        .IN5(n1444), .Q(n1443) );
  AO221X1 U1971 ( .IN1(n359), .IN2(IFID_A[8]), .IN3(n358), .IN4(IFID_A[7]), 
        .IN5(n1445), .Q(n1444) );
  OA221X1 U1972 ( .IN1(n358), .IN2(IFID_A[7]), .IN3(n357), .IN4(IFID_A[6]), 
        .IN5(n1446), .Q(n1445) );
  AO221X1 U1973 ( .IN1(n357), .IN2(IFID_A[6]), .IN3(n356), .IN4(IFID_A[5]), 
        .IN5(n1447), .Q(n1446) );
  OA221X1 U1974 ( .IN1(n356), .IN2(IFID_A[5]), .IN3(n355), .IN4(IFID_A[4]), 
        .IN5(n1448), .Q(n1447) );
  AO221X1 U1975 ( .IN1(n355), .IN2(IFID_A[4]), .IN3(n354), .IN4(IFID_A[3]), 
        .IN5(n1449), .Q(n1448) );
  OA222X1 U1976 ( .IN1(n354), .IN2(IFID_A[3]), .IN3(n353), .IN4(n1450), .IN5(
        n1451), .IN6(IFID_A[2]), .Q(n1449) );
  INVX0 U1977 ( .INP(n1452), .ZN(n1451) );
  NOR2X0 U1978 ( .IN1(n317), .IN2(n1452), .QN(n1450) );
  AO22X1 U1979 ( .IN1(n1453), .IN2(n316), .IN3(n1454), .IN4(IFID_B[1]), .Q(
        n1452) );
  OR2X1 U1980 ( .IN1(n316), .IN2(n1453), .Q(n1454) );
  NOR2X0 U1981 ( .IN1(IFID_A[0]), .IN2(n351), .QN(n1453) );
  NAND2X0 U1982 ( .IN1(n345), .IN2(IFID_B[30]), .QN(n1419) );
  NAND3X0 U1983 ( .IN1(n1485), .IN2(IFID_B[31]), .IN3(n1422), .QN(n1417) );
  INVX0 U1984 ( .INP(n1455), .ZN(n1422) );
  NAND4X0 U1985 ( .IN1(n1275), .IN2(n1456), .IN3(n1455), .IN4(n1457), .QN(
        n1412) );
  NAND3X0 U1986 ( .IN1(n1486), .IN2(n1003), .IN3(n1487), .QN(n1455) );
  MUX21X1 U1987 ( .IN1(n1458), .IN2(n1459), .S(IFID_B[0]), .Q(n1415) );
  AOI21X1 U1988 ( .IN1(IFID_A[0]), .IN2(n1274), .IN3(n1008), .QN(n1459) );
  INVX0 U1989 ( .INP(n1456), .ZN(n1274) );
  OR2X1 U1990 ( .IN1(IFID_A[0]), .IN2(n1275), .Q(n1458) );
  NAND4X0 U1991 ( .IN1(n1488), .IN2(n1487), .IN3(n1005), .IN4(n1002), .QN(
        n1275) );
  NAND2X0 U1992 ( .IN1(N223), .IN2(n1269), .QN(n1414) );
  NAND2X0 U1993 ( .IN1(n1011), .IN2(IFID_A[0]), .QN(n1413) );
  NAND3X0 U1994 ( .IN1(n1001), .IN2(n1005), .IN3(n1003), .QN(n1456) );
  MUX21X1 U1995 ( .IN1(\regfile[0][0] ), .IN2(AluOut[0]), .S(n1276), .Q(n398)
         );
  AND2X1 U1996 ( .IN1(n1460), .IN2(n1461), .Q(n1276) );
  MUX21X1 U1997 ( .IN1(\regfile[1][0] ), .IN2(AluOut[0]), .S(n1277), .Q(n397)
         );
  AND2X1 U1998 ( .IN1(n1462), .IN2(n1461), .Q(n1277) );
  MUX21X1 U1999 ( .IN1(\regfile[2][0] ), .IN2(AluOut[0]), .S(n1278), .Q(n396)
         );
  AND2X1 U2000 ( .IN1(n1463), .IN2(n1460), .Q(n1278) );
  MUX21X1 U2001 ( .IN1(\regfile[3][0] ), .IN2(AluOut[0]), .S(n1279), .Q(n395)
         );
  AND2X1 U2002 ( .IN1(n1463), .IN2(n1462), .Q(n1279) );
  MUX21X1 U2003 ( .IN1(\regfile[4][0] ), .IN2(AluOut[0]), .S(n1280), .Q(n394)
         );
  AND2X1 U2004 ( .IN1(n1464), .IN2(n1461), .Q(n1280) );
  MUX21X1 U2005 ( .IN1(\regfile[5][0] ), .IN2(AluOut[0]), .S(n1281), .Q(n393)
         );
  AND2X1 U2006 ( .IN1(n1465), .IN2(n1461), .Q(n1281) );
  NOR2X0 U2007 ( .IN1(n1491), .IN2(n1492), .QN(n1461) );
  MUX21X1 U2008 ( .IN1(\regfile[6][0] ), .IN2(AluOut[0]), .S(n1282), .Q(n392)
         );
  AND2X1 U2009 ( .IN1(n1464), .IN2(n1463), .Q(n1282) );
  MUX21X1 U2010 ( .IN1(\regfile[7][0] ), .IN2(AluOut[0]), .S(n1283), .Q(n391)
         );
  AND2X1 U2011 ( .IN1(n1465), .IN2(n1463), .Q(n1283) );
  NOR2X0 U2012 ( .IN1(n1006), .IN2(n1491), .QN(n1463) );
  MUX21X1 U2013 ( .IN1(\regfile[8][0] ), .IN2(AluOut[0]), .S(n1284), .Q(n390)
         );
  AND2X1 U2014 ( .IN1(n1466), .IN2(n1460), .Q(n1284) );
  MUX21X1 U2015 ( .IN1(\regfile[9][0] ), .IN2(AluOut[0]), .S(n1285), .Q(n389)
         );
  AND2X1 U2016 ( .IN1(n1466), .IN2(n1462), .Q(n1285) );
  MUX21X1 U2017 ( .IN1(\regfile[10][0] ), .IN2(AluOut[0]), .S(n1286), .Q(n388)
         );
  AND2X1 U2018 ( .IN1(n1467), .IN2(n1460), .Q(n1286) );
  NOR2X0 U2019 ( .IN1(n1489), .IN2(n1490), .QN(n1460) );
  MUX21X1 U2020 ( .IN1(\regfile[11][0] ), .IN2(AluOut[0]), .S(n1287), .Q(n387)
         );
  AND2X1 U2021 ( .IN1(n1467), .IN2(n1462), .Q(n1287) );
  NOR2X0 U2022 ( .IN1(n1007), .IN2(n1489), .QN(n1462) );
  MUX21X1 U2023 ( .IN1(\regfile[12][0] ), .IN2(AluOut[0]), .S(n1288), .Q(n386)
         );
  AND2X1 U2024 ( .IN1(n1466), .IN2(n1464), .Q(n1288) );
  MUX21X1 U2025 ( .IN1(\regfile[13][0] ), .IN2(AluOut[0]), .S(n1289), .Q(n385)
         );
  AND2X1 U2026 ( .IN1(n1466), .IN2(n1465), .Q(n1289) );
  AND2X1 U2027 ( .IN1(n1491), .IN2(n1006), .Q(n1466) );
  MUX21X1 U2028 ( .IN1(\regfile[14][0] ), .IN2(AluOut[0]), .S(n1290), .Q(n384)
         );
  AND2X1 U2029 ( .IN1(n1467), .IN2(n1464), .Q(n1290) );
  AND2X1 U2030 ( .IN1(n1489), .IN2(n1007), .Q(n1464) );
  MUX21X1 U2031 ( .IN1(\regfile[15][0] ), .IN2(AluOut[0]), .S(n1291), .Q(n383)
         );
  AND2X1 U2032 ( .IN1(n1467), .IN2(n1465), .Q(n1291) );
  AND2X1 U2033 ( .IN1(n1489), .IN2(n1490), .Q(n1465) );
  AND2X1 U2034 ( .IN1(n1491), .IN2(n1492), .Q(n1467) );
  AND2X1 U2035 ( .IN1(n1468), .IN2(n1469), .Q(Zero) );
  NOR4X0 U2036 ( .IN1(n1470), .IN2(n1471), .IN3(n1472), .IN4(n1473), .QN(n1469) );
  NAND4X0 U2037 ( .IN1(n294), .IN2(n293), .IN3(n292), .IN4(n291), .QN(n1473)
         );
  NAND4X0 U2038 ( .IN1(n290), .IN2(n289), .IN3(n288), .IN4(n287), .QN(n1472)
         );
  NAND4X0 U2039 ( .IN1(n286), .IN2(n285), .IN3(n284), .IN4(n283), .QN(n1471)
         );
  NAND4X0 U2040 ( .IN1(n282), .IN2(n281), .IN3(n280), .IN4(n279), .QN(n1470)
         );
  NOR4X0 U2041 ( .IN1(n1474), .IN2(n1475), .IN3(n1476), .IN4(n1477), .QN(n1468) );
  NAND4X0 U2042 ( .IN1(n314), .IN2(n309), .IN3(n308), .IN4(n307), .QN(n1477)
         );
  NAND4X0 U2043 ( .IN1(n306), .IN2(n305), .IN3(n304), .IN4(n303), .QN(n1476)
         );
  NAND4X0 U2044 ( .IN1(n302), .IN2(n301), .IN3(n300), .IN4(n299), .QN(n1475)
         );
  NAND4X0 U2045 ( .IN1(n298), .IN2(n297), .IN3(n296), .IN4(n295), .QN(n1474)
         );
  MUX21X1 U2046 ( .IN1(n1478), .IN2(n1479), .S(N254), .Q(N324) );
  OAI21X1 U2047 ( .IN1(n1480), .IN2(n1481), .IN3(n1482), .QN(n1479) );
  NAND3X0 U2048 ( .IN1(n1483), .IN2(n1001), .IN3(n1269), .QN(n1482) );
  INVX0 U2049 ( .INP(n1457), .ZN(n1269) );
  INVX0 U2050 ( .INP(n1494), .ZN(n1481) );
  OA21X1 U2051 ( .IN1(n382), .IN2(IFID_A[31]), .IN3(n1483), .Q(n1480) );
  AO22X1 U2052 ( .IN1(n1493), .IN2(n1001), .IN3(n1484), .IN4(n1494), .Q(n1478)
         );
  NOR2X0 U2053 ( .IN1(n346), .IN2(IFID_B[31]), .QN(n1484) );
  NOR2X0 U2054 ( .IN1(n1483), .IN2(n1457), .QN(n1493) );
  NAND3X0 U2055 ( .IN1(n1003), .IN2(n1002), .IN3(n1486), .QN(n1457) );
  INVX0 U2056 ( .INP(N255), .ZN(n1483) );
endmodule

